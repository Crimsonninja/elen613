







module uart_top(wb_clk_i, wb_rst_i, wb_adr_i, wb_dat_i, wb_dat_o, wb_we_i,
	wb_stb_i, wb_cyc_i, wb_ack_o, wb_sel_i, int_o, stx_pad_o, srx_pad_i,
	rts_pad_o, cts_pad_i, dtr_pad_o, dsr_pad_i, ri_pad_i, dcd_pad_i);
	parameter		uart_data_width	= 32;
	parameter		uart_addr_width	= 5;
	input			wb_clk_i;
	input			wb_rst_i;
	input			wb_we_i;
	input			wb_stb_i;
	input			wb_cyc_i;
	output			wb_ack_o;
	output			int_o;
	input			srx_pad_i;
	input			cts_pad_i;
	input			dsr_pad_i;
	input			ri_pad_i;
	input			dcd_pad_i;
	output			stx_pad_o;
	output			rts_pad_o;
	output			dtr_pad_o;
	input	[(uart_addr_width - 1):0]
				wb_adr_i;
	input	[(uart_data_width - 1):0]
				wb_dat_i;
	output	[(uart_data_width - 1):0]
				wb_dat_o;

	wire	[7:0]		wb_dat8_i;
	wire	[7:0]		wb_dat8_o;
	wire	[31:0]		wb_dat32_o;
	input	[3:0]		wb_sel_i;
	wire	[(uart_addr_width - 1):0]
				wb_adr_int;
	wire			we_o;
	wire			re_o;
	wire	[3:0]		ier;
	wire	[3:0]		iir;
	wire	[1:0]		fcr;
	wire	[4:0]		mcr;
	wire	[7:0]		lcr;
	wire	[7:0]		msr;
	wire	[7:0]		lsr;
	wire	[(8 - 1):0]	rf_count;
	wire	[(8 - 1):0]	tf_count;
	wire	[2:0]		tstate;
	wire	[3:0]		rstate;
	uart_wb wb_interface(
		.clk				(wb_clk_i), 
		.wb_rst_i			(wb_rst_i), 
		.wb_dat_i			(wb_dat_i), 
		.wb_dat_o			(wb_dat_o), 
		.wb_dat8_i			(wb_dat8_i), 
		.wb_dat8_o			(wb_dat8_o), 
		.wb_sel_i			(wb_sel_i), 
		.wb_dat32_o			(wb_dat32_o), 
		.wb_we_i			(wb_we_i), 
		.wb_stb_i			(wb_stb_i), 
		.wb_cyc_i			(wb_cyc_i), 
		.wb_ack_o			(wb_ack_o), 
		.wb_adr_i			(wb_adr_i), 
		.wb_adr_int			(wb_adr_int), 
		.we_o				(we_o), 
		.re_o				(re_o));
	uart_regs regs(
		.clk				(wb_clk_i), 
		.wb_rst_i			(wb_rst_i), 
		.wb_addr_i			(wb_adr_int), 
		.wb_dat_i			(wb_dat8_i), 
		.wb_dat_o			(wb_dat8_o), 
		.wb_we_i			(we_o), 
		.wb_re_i			(re_o), 
		.modem_inputs			({cts_pad_i, dsr_pad_i,
		ri_pad_i, dcd_pad_i}), 
		.stx_pad_o			(stx_pad_o), 
		.srx_pad_i			(srx_pad_i), 
		.ier				(ier), 
		.iir				(iir), 
		.fcr				(fcr), 
		.mcr				(mcr), 
		.lcr				(lcr), 
		.msr				(msr), 
		.lsr				(lsr), 
		.rf_count			(rf_count), 
		.tf_count			(tf_count), 
		.tstate				(tstate), 
		.rstate				(rstate), 
		.rts_pad_o			(rts_pad_o), 
		.dtr_pad_o			(dtr_pad_o), 
		.int_o				(int_o));
	uart_debug_if dbg(
		.wb_dat32_o			(wb_dat32_o[31:0]), 
		.wb_adr_i			(wb_adr_int[(5 - 1):0]), 
		.ier				(ier[3:0]), 
		.iir				(iir[3:0]), 
		.fcr				(fcr[1:0]), 
		.mcr				(mcr[4:0]), 
		.lcr				(lcr[7:0]), 
		.msr				(msr[7:0]), 
		.lsr				(lsr[7:0]), 
		.rf_count			(rf_count[(8 - 1):0]), 
		.tf_count			(tf_count[(8 - 1):0]), 
		.tstate				(tstate[2:0]), 
		.rstate				(rstate[3:0]));

	initial begin
	  $display(
		  "(%m) UART INFO: Data bus width is 32. Debug Interface present.\n"
		  );
	  $display("(%m) UART INFO: Doesn't have baudrate output\n");
	end
endmodule

`protected
b8dN.;:PN^6b]R^T60a.9J3<)U&ObGXNH,eJ3=DLE[<J._)@C7SH()/LBL6D\QWO
cedB?Yb(1(8+.&c.K68g3ec(I&EdP#NFP\+6D^S^+0(P0EPNILg)WWZLdPDaGUNV
JC6\1gc1=]FSQZZ:]#/:fJ52&=E16]8Y=<:3<KC=YbZa<RTFTOX8L1S40/\?RH53
Y0LfU7^I(f667_HZ:.\.,-3I=:,?=:b_=aNdMBc#+W#)&LJSWN[STBF8ZWB82Q@d
97X9TG(&:12ZS7SWVaBV1UUMLa9+f/A<PBg80@Rf^+7U[WT40+.QDN5121[f2JN_
b]&MbO-V>R1#NV],KMMaTgEfTMQQN2F8L6Mf3dbN_Z,PC_^BaAV@^dM-?A,U@dE=
M<BU<<U7gH10MKHb:WESN&AfC5@>F<eZ]e9WBTXg2+,SZJX=5A/OdM/X/Z6TbIDW
,bXRJH9_LF8aa:22?65^.1>U<F?1,#^F5TC<Z2PWR>7,.(2PVGfDT6Q7]@DGX9V)
IU50J3]\8FIGE2GN2[CMgW#a?^;3d7#&.AZ#SU0(?W)[aV3DGJ9eO4,Sf[Z1MIdP
,Yc--G-5];Y,d/R=dYc>fd73Se8e,47VW-D,3.)H;4(d9;H@cQ\LNCgSBME6U_FB
DO+5>Y+JOg#+-KC_IKH\^-3S2(g1U#O/+4/\L?XK,VG?BWW+U#TF]0:g:Ob)N3gX
,cP&@;GbZ_R9N54N.TB8PWdeGDASI9)-=0aTb6([OdNb23FfJe^[a9#+=f-b;c\(
Q#13(HCGaLfJWS_^Ad\R@;05KK_UHH1,=@55)Q>,d29\T\0P-+/>5P=3\YBS<DgH
_)?ROe<;]N:HOb[WA48(C2EM6HEcESU^)W>eY4&\&2PMNEAI<@FJGE:RV[Z^8)>S
KeCLddRg^=[DU7[A;cC5==1V1#:888R=9B&_D&HF>8+.a6\<XD]46SI1IV(L)WV1
?9UD0HgWX<[cBGd)Y>=(/9@WZ[A7+-QB&89(F&UTcV>]_@.L\0dN;^eJ5N(-8Rc4
CEdPTe3c_-e0fI.)_O(NU[T;Ia0B\J<1>IY58W:<#\=eL]001YeM/Dg1Z7]Eb,_O
Y^f2)fJ,9JH86=)Z6@:YT(&<7CCdYMV-7X7W5#AW-86HEOWe?C+:P]-]@f24?56+
Tg9(-M(&;/_9DAR8a@ZLe1=8TdOOS-O8C=-FV50M=^Y5_U.K_:OX[4;>@Y1P,+PT
KXN3^R5QGDRI?Y^RfWfQL12BZeVP05CYU^/H(G([caBe5DS7#d;EQ6OEf(G(D?cM
;C95;H9ePc0N;HB7IcWNg[V+cS4PH.+=<0Lc-U6Q\JZ0ba.B:_[,(H=(d/=0LR90
I2UO[dC?8[2VFKMM?;]4@b1YQ8G&Z/5aBM/[44Q)/C4/M^N[B<:3a/Wd_dU(7#@/
WWfCR@&OLR>G<+Fd10^4^20V&DGO1PdMWW.01Eb)<Z\C)[_3B&^QTY^7]6.PNMVS
L@>_;]&?>K_YgQR4&b46g)X[V)YfU++95gKEDdXR#XK,IMV^8Ta9b,8Z_TH^=RQ+
&O7E5I,[JQX1ZG^U<N6/?YZ/Bdb\gPgPMFaFU-<(a2AJ<;?Mc;6<07aOJTdL@K)b
^AEOD4OIA]G#6GJe1Z29UXF5GTVJ1/)(HY_FYdCb#b=1EP/(F-0J>.-XH;Tfa?@W
IgL3.TT?\Ya.]\<LIFf&+AZb.SAERc+QM_T;&K@_)_M2G?-Va=>_:Q<=[G0>1=D)
/1E&_W=^&J=-EG/ePU#ZXY096aeVMEI]&9X\WBFQ+YV/:d)MRFXC4ER#a;)8CbfJ
X>_^>_8Cc?&:ebW2VBbWeU1c7g:Y7?H1Y\PG:BQX>^4S[UW&4aM?U1(WM.)3?a3M
K?JVNY0B8.EJFUI<+M21_3G/L)@06M>b@O3<]=f,e6L+aa3LdSQ#\[/6abO/.VH<
XcYKN]Ad>)<NTJGHOTP\+RH.L-=,0,GTXf6LObMEHWB/5ad^Sc83WEHB:-\U:RZC
G[A>9U(2fJFgW11R[#S@1Y].7(db;L.0;FB+XVSg<Z<eR4]V].NRa2WOY7?;g8Pa
Jf1SD[8M?IA.Wd<SH9Z,TD1gBa]9MQBf<,1G]S4e:5[\Zg-[KRg5_<G4)Aa;TMV#
Me/CL.=b&0H0IeO([gf<A4JLFS[-=3U>f][eTSB4)<-CGAH#\=<.4Z4aOc10->>8
BT&E8E]fQ\QBFH3T.N9gI+c4B[O031D:I,>]PX[Q2U+cEI3O&W@VNd:c;UJLGAYd
ccN,&TIfcE+e_@eELg=(&[R53&32P(XJ_d;S(YI+4OO?0aSN1CIJ51PJL5L#26X<
b7W?P7O_2.a8Q5[PHN-2daXcNU:CRXKNK^RAIMH90)OIZB0)=5gQPI35-YgaLQH<
bXL:UI\HdUE-&Ib62D-;&>+U3gATVcYgLaH8X?g.A,AO34NF\(b+E+^YM/\6Yd^>
VbcB^MaCVb@[OgfO=_?-M/MdSQ=gaA:JEZ4C>]de@CfCKILVcL@:>^,Q_PN?,aHV
;.EJ.fMF5aIJ&>RCc/W?:E,RW88bXKW9;;c-EGc-Ob3[c.c6fC<NU2P<DU5FbF7E
ed4VTJQb5cGQOe[>/QFNJKEIF3VHKb)I[;Sg475,8W0Q)7+B;+cNKJ/?D[P1)&;Y
ZY_PEIQP4\&YSJ.d_EU<fBFM9UQYBVWY47DG,3CS&GOCP];G,.;+CaF4dP>Gd;J-
G>?.(,Jf>K(RZ37(Rd:KHa.3TQI),=_V(&FaeFAL24Y2/g&NX2:@&Rb60NR-XB#O
+3VEN46T;4ZgL/f,dQ[KQfVAJN_c+Z?(,WH;0#.A&)B3KJ1QYUg\8LD7I,VZ&=TM
YXDbESEBH9cMD38QQ<;/0aK#M-^>e/.H#@?bJD-Y)E3#Y84+6AEIZa<OW7,V>QZ?
2I-PYD])O7_XZYgJ4#3YRST1L+GSKX@?.CEAf;@CfeGJNY4X?5#[D\[YH&=N8\>)
K\)TN0f@<+1-gfYQe7.66MS5.PWIT@H8YPLVV_ca&(N<3.G3Xc=@(.UL)H;7?cQP
4?UEc6fMc@V;C8aQ)cA)&PUX>[O4?H@aYK;2)^-F]NV@Q,)FLf5<B+))6^\D;O14
3+?d\,W:1XI4/(D//;S0J[\bH.IP?J5WC&R@b)MJW4?ID_b\/O0_HM,8b89Q.+Gb
&9LF]ga_NZ+YcM/M_GLe>NS,S+0Ag0AdCe^&+X_Mb^)MZH<5g]NC2G.UX.EIRB-d
YT?Z,?M,O-TReeYC\\/(40K7Q=O07?Wf7V=&a)SU1TZS?b9O5NIU0cUH-J^JO8FJ
<JG-Q:A^>BLRGF@4<aeVQ2Q-[Fb:,?O1?OT_Z+P3?Y(Ja^_81JJM<:SH=#^c.I9_
T;DP\BNTHY/XK]]Y[d.\aS-:?bbYS47/3:3,QUN_F@F.afWg,CFWE73X>4<#:E=Q
60d</E3AEaSeP[eSa[38VH9(^:?]O44K-S.CgVTGW+(&d=Q,<GHR/]R7X@09O:=I
13<0@QYTeX=KRNcE;_2dBg_6a^MI->LCe],9Y2F?e#BSFFL[DO/>]a8XVdb8#D)&
:LV1W\:D&-,7QfLA;BO>ZW@[XcR:7fccC^KSaGLQF?=M=4Q-PEd0DEKB#X<8RH20
J5E/KIBQab]L&E5-IC&U7&R?O2\5#OE=O&J9SEX(&#U72<U:JHQ=64/:D#)ce-fK
>[USTWVeHC\SSB0^\KIDP#(X_W#Ie6B0&W[Be2V5Zg(#9P3/F^O,I[B7ERZ8f#2c
deG@[D&35)a+#,+?Ce>/,#E]9-dQQ\GIdPF^B6a.]-8+Y;a=\B.,\>ff-SE#dZR?
gRSLPC_P39PM)MQOTOdf0b+L@1F(/>>>aP([Q^63YS(HOK@<Md+R#U2J=fS<_?cS
a<^@f3_Q:/PM[<V/XNbGHPd]Y:1\P.Nf.OO7PGWWJTTFZB-?C:09_6dX^:RJW#[,
YEU,M&e+Z+?M+>U+R2P?GK_8EJN\<DAVLg@;B;KSMUa@&\70+J3J\/V;EQe2/GUd
I5b1MI5(6,:BW1MT:EV518[[N/I5O:\)5eXXEg>f+ST7ff,_Zff_PEa1O()5)X.P
>>^DYA=>d7F_fEOcKP#TVPM5SgO+3JBS]:K&<BI?d((<6FP?e8CF@(Tg^.,X1CQf
7LMXO[d<^e1/E.,)(X=D+434Z5PWW(&CUH1IY/BZXCEEDa0IPV?,I#;a;V^bTg@Z
.-GFVDI^DT\g2348NWP+fA.KR&ASHJbU4XB@R(ef,)L.7#.+fO[BE_./BPVgLD<#
PK1\]3=<<]7S5?33(#0:CI]V_O3feR4H30PJ;8:S]gcSU#\@T[#A-NI#L^e)3ZOX
Jg@),;)4c1T?E[D=<9MGL:a6#]CJBX]HH6@RS;8b^0<[DB:.N83C\<Q^Q5/@AaAW
OR<cTYB._cda&/X9>_,U:./^GTAe#^dSD&(5TM#PS[XaBEQ&cS,+^FF1fbcVRD6_
3@P.87=..0D3W/WR6+S1Qf,W)2Zg0f0CbP=1V@A5R;Z&_LZ[[bU^V3R8e[PY-CS3
=^2TI]W)XT)@NO0XUc@FU?5QUY6Ze52,C]UdC>TR@bIfD_/:_=FLO.FRNF[<SR+R
;;,ARa]J&S6AKZfF3gP6O?/^W7CWIZ6?K-NKO=FT0H(e;-\#fI979H-14I)6+A\8
MHQGBEcaVgL>JU-X7-^?KGbDI\d].,,^4CdfEOUB2E8eY,J;)>7aF#J#O&T^_^A1
FWX@MLR.0CB>3db#=:;Wa:S1/#>WVUX/+]K\)M0=).,VC7B^MWD4-V_V]=DIMQD5
BNR:LY(DObZ=AHabc?[X[A8VF3cM<MM4?8Q^H)N6(LWVYF^BT^J5E&1EF5D3U)/9
-T=L&4+:TgTNOfLSL^EXF0DIL=a?1ZVbFN:B8+dF+#XGf#W@LT,>+9\KL1;Qcb8E
2:0JdT^JX=_cG@&eE&#LS].e,Wb0Uc:dE&-GX[86Y;G3;09FLFUGLUYgUfTS3ZLd
B1P)cT/RSfScWDXP5HDPU56I6cHL^@GFUB-7(C@<SZF>Gc[2?Z6cP];U?RCJ=I\&
=SW.U)ZMDHI+@9\7><Y1[HcC7b-/[/Ig9XRW+(+T&A/UDNYU_<NWW6)YH7?_UUD3
C3[X4ddZO6W8AUUF^U@U,?UX<Y</eE^\]PBCbS2\2T.DVYPR1[N3fJ_<.f[5(O,U
KX[G;1.5=:CGfDQ2QdDd^I2@Ea(:b:b(FEN())_dcU&+-L((]Te0T3#;T[FP-R;8
7CNWO;.7B0<9>\74T7P](KH7cC=.:3UaVTN_TXWb5g/dJS0T41(HC.8JS@@?8\MF
VS3-=gab^[ZaS2-^gDa;4QM#aa8,#;?Sa5JK,1=0X1f)U9P,7PBXSZCD(1>A0g2.
<I4AY4CB363>&))RI[I7PPKC8R4VS^aNFLBT)O]Q#+4R@/@?FE125U/AT#5@5JD3
\K<(K6(13UdISB)5c<cBUZ]ZV(A7S1H-KW2\(-G)@?ALC2XKDEN)S[1@EER.e]YD
FYJcAYOFD\^X>F,/A4U_O1^K>Z7@R?dKI@fC,J>;M(5\c7Jc@7,P3A)=?>f:Bg5E
Zc8FbG1,X;KdY_BRcS(SN/Z,2?:9_P3eTC-Jc_LF?V,OVb59?KZWd]FeIc<RVIa6
;-IBLV4]6]L#Uc34ED?8I^=Y<&cLL4F1Z9&>1fBMeDSNQF:GJAF(-6bI);&_OOaU
-\]DAR9\33TCS#c#)MAH>+7_:^7G\U6?)#Lb1Z^\;+<H-J[8cFATBdV(fg-U@?OW
:VF=^d8EeNH\]ZB:X\#L[V]BH6c/6-&Z:Ug.?69.F9E-)(3WTETI+ROg)(92?+GN
^O_a;\5OLZTB)F?g1C#XHEL[?;R<WAV/NdI9?X6\),Y:9]@V#W6=cZ-_^-=ECed]
QO:4D8.UZ_,6I.1dP(N8fb>)fF9b+][.aWA<0RaCc3KJ@KfLF#)/&AdL4bPd5=dY
@EX)>PX7ITL1>UUd>A?C)?E/E&K)d][#+O-ZI25#^1fKWD+\8;XU=4^JO1CAcU_.
cb<R10OD^bM+;4g?D#gE+CCNPA\M/[?Sc0T9]L2,/Z98PFDAKOMLEHCWZ]Mc5S>[
=dgE(OB.NMLM?+NW:T#OY>gVK9>_GZ1&(QUR>9(\HY4_3b-3G^6MGUJOa(0YQA+F
:bF#\@fa/DObBI_<&Cd;aKA-;_2+c^P/4;c5eX))X6?1G]B3^GT&6)&HFgP[LF^Y
d^BDd+O&\@PH7+?YB_[T#\bZHWT62-VG8IM3@@d&WdJANb,7aJ#L^-E[JG+;1bE#
QCJ&]g=M[>&Y<DggI4ZTUAHGXE-e0A#NAN]HZ+(E7?EJ(#ge1\_=#^RfA8PXV,8H
QTC&0XHQebN5+2C[a_D8SgDbC1Ue2XCbgYP:Sc6OFI;L/>7?R]##=(AIH.2JS;P6
dF/8KU&>4(bE<FNd<(J=W(,T>>X/8..:B&KX)^3LF#F(@+Xf,LO@MY0;7#<W.\&=
+dJ7I7@SPQ)ZcWXI,5]S3EOQVBBNTRG)C843^RdT+FNB<_P+BUH>]QR(E+](?]R(
T(UL9:1?&G]ZOF8MLR4?F)8&K;[E6daBf]0L\Q^+CXe2g^5^,MFAS#d9SXdBGPMT
b_/Sa,SDN=GQ7[-28GFE+<1-6c#A8IKLZL@7H7gdf]?)\2gS=^GK#J.G2K-.f2&K
<SEBYHZM3)7&3D:fVYU.fOB&NQFW)aW/W,dO&9f.>E;M4d2^(;/J,BfA<S?:c&3>
)2W/?,(SDeQC)Q(+-9=7+R)3L,ZE5>DcF;YN9FFMb565FX;<U_.:eY/\6M^=VY=P
TLZ3TVB6Wd;32#_DF^38ZI+DHK=SQ0O0V\C1/-AQ,XNDMXJ;3183OT]X+fUd;dN8
217I^4(S=:N-10@9;fGDa(\7UGXOdPQ[^dD?JK3Ugf=L+e:SC^X;MRV;5=(d_M)I
NU=IGH.7\_e;<EV-/LW<(7A81+L9T4a,56fM\P5OVC,>Df,,KYdg(PYed/&#VZe2
-Q/FI.eea.R=X#/DP5gg(f]\OgfE/3d(XcL;/_,80^cBRM80M;]<,B-C\JQ7dLW;
BY7=\=XR]/.?,XICD/U/H)5-?,Fc(DUO?\0a(M5Da3S(.<<@DN&V>S[(Y00aS8aD
1<(A>U]74#(##H5S)7f^Pd.MRJLPZA\B?\&SR0O7d>1?Vf4NH/VgQ<TS+5&bfE_W
<0QQg6C;#BcBaE6WX;.WYf/1VD?MHHR8]\(D,7+KD[]3)\<P5Ic6A?PK/)K_K^8U
6g<,K:f=/=NM?BS^QMUg0c>A\NVPYI3f;K]cYU_E<A7[Df4d;EHK[b[HDWCJX>A/
>a]gf_KAJc,Q;d;VK82^+Y)32Y[E4eVXfdB:LL>W#T_]E9eE7WA8/>c+5)+/MC07
0IM8COQ89a^Ub9<aM(dRdcGPRWZ-eABL0/=,=#GUOOV>bK(APL^;MRU6.#;_[[/5
R92D+B--/[f7Z^V#QGOBRN\58e4MgHOWYIa8NOXgf9cUgJ\G\(885Q(K\g@5?:Na
4L^#eY]#;8b7<L=Ce55QR5R729>Q-G[1R,5UE]CY77)2I7?7EfAfEB>2:d&[O6>I
ZB8&X)4<:IUBV&4beSg7<O=YCKafTCOBRQU7cU:41,cW;+W/FYWSXTT311@]JC,L
^&0:N>e5W8Q9e)U,<[&AD0M7cQ#I5Wd0RR0>:971f+,Q8,230GWf>&H1.)8NO,M3
&2J)2X236CA2A=4[:23.f#A3\&1EZS#52-^7KEXYFb[1)-1AH94&U,@SOd)#]7O1
S^&T]Q0;e/4/]VUHO.^ZB]bJA^dg=-c_FN96SQD&4D>J=E2[O;@P-\LHC4Tc;AgS
<<,^@UYPB82R-]cKHV@8@E9OIb@-YRWa?]M<g#GdPe:M0b<)5]SAbWBXYf#>.0/<
FPd3(=e==H>6IQ)K3&_@0-\^_YM8HeG7]-S@J=I9>]Jc;?PacfF<VgD7Kc(eZFY=
^JHA[:#(P@AP3WI9?H3[_RKT+C\GW:e[7)<09BKY0X1caegD[B9)FCBdSJC4\X:5
UV#DQ#_>V[bM&\(I\FXYbB6^5=317@aCJ9@gEgK4QH4<HJI@c;S,;3X+a,0d@O\F
\^7Xa]#P\98]0UfRZcD45,Y8.QfIC[FZeSQ;1>;+aaT:I,RRH9gd_0T+X?]G<:JY
L_f)[8.J0)A\Cf@K04FA6d1Ab3A82@VY4a6)9\QeO(0K\QP^#]PN-&1H?-SXB@Q4
MGRA(X(a6)eNe(b_NVfA/M+<4b?#FQLY2d0Z3g)-;ADcbAWV[O,@:;Z1e4;c3T?d
BbdLaF@](ae<MBW??f(^Y4Abc@BQH7JJ\)7],<V).>UVB#WgK]0X\geQY)fOR0aN
+dDWJ4MIE65QO18<>#U,+1F-6TYgPAC:=#6>-&>IcR]\b538EL&c_=:M&aX)E(/8
2C@TWcg3C4:V4PBc]<VV@+UF@0.Q2;#EV5?F=Q4e-XFE-6Z:,I_;)_O(TOg3-FQ0
&O5Ba3>57:cZc=d_a9I/QgfW,ZDBJEB)3cc#:bV9NQa:Cg#..N5]2a7=4:G>gWa?
e+=A<?c.d4OHW,b.]@Tb5/EN34WaR.-&b&TO(&+f=0C<g[XHY7a1Xd)O-HJcF=^9
G@21)\8_Z_)LJYC5G5XK,ZYC2^[2S:HRg55Qg-,[XU36F+VGX64a=SJR66,B^YF;
#8_]WM.^>5=]>6:Mfd]T1WCeNZO2d,RH4dc1H-/U<Mf/J-]^UET05^X7&2F#8NL2
F=ENA258C/6Q&g3]]Q]HCAW(BKe+0&PN0V=73374&9g97UC;Q=c5?dVO^0AcZe+O
9>bT-8g+f++/#bf+F8>S=L@gKgIeC/XV^R)GK<MT]JJ@W7S=L8DcbV6IbNVHbY@P
4YKW8-3e_&M786:YC_e@=L^)/U)?+bC4gH0LJfTb597XP<U^M8&\39U=c,.18=VY
W&O<7\#bCY:U9_Lg(O4(03/-FTG4d;5=QZD:,N2OPNcJH^_N>IH/aFZgO0CB=5Q2
C]IfBYN5fT@+g3:Q2?a?[8Y(K4[d2RAM>IM5X066-Q3-9(1,9#MFM9gN,V[T6[B\
#X&ZVEE@5JVg>dTZZG,4,T-b(154e55R_O7UIUK7U@0C@:FLWNXR7d/-Fc./<d@]
dB1\_FSR2)T_Q5e5-a_RPbP66Y\9g<CNEYE#eIHY?C/^U+DDME_>7_:IR\<:NXE>
17@AO=8ZOd2Jg&:cVcNY)/7ZA3Q1+bN\+R8J,G#bEI<\O;@cS0RgOe3ZR&GJA>/P
VLTa+<UVGA:;Y;K[CC:f6/TFf(KL,1b2a1__8cHAH>S7]CIDdJEWO:8ed(bU6\2,
UeDJ\80GS947BH23/IJO\3DECT5>Tdb].@QJ04#NKc^6VUXC863\cPfH+F8AERD,
KV(EfMOS47G@(TQaZ@2F+(6[P:@^ODY.-bJ)B+#(Kg.(N/\SZH&cYWS^87V;^+/5
8,)F>LgR4<;&WfTf(f4aE3@\D0>A>gV(2T;0-I\<>VRa2S=45Y50@,9T[)f5)\e-
RH@+0CKO8EM48)ea1\TQ/N6&d3G#JLX@fCaUH4Nd:,5]eN;]N:++]c-8P_/R<;8(
-&^^^TV,G\<c4VD<)556]L9:da=eSJD=IN7\IDSZ:^S\V),>E2KIeNXX(O=CLS3g
I5DN<\fd?cgC1#7I\3&AYPW&[>bLU^6X7X<R?LP^&RfW.\a5:9N?g01,#BM;&3E<
(PQbI3[B;JH#8a=C?(M(_QE:<20WTC+_LSS)HXA1/,1O]MP,M/fATRKPAGV7AT5Q
bLI_b(:6<Df#E3U8@HJI6-1[QABb[85N0:POO-C,#BF(a=9X>37D,fZ3G>_=M5)^
9X21Q8^/5_,+<AQ79DCX3GLOG/&X:8O[QK<1C2,B?OONK8G2>Z&+>0df.L^+L7_;
Kea4^fgI/VP5)04O\A]@NGH_;V34e9I9)M8WPYfY@1Z3RL2^KZ5eCHU;:4T6]#G^
[RKN/19[+3_@,F30R_(86T.F(fXI2T4gRQX-\W_2=M(c,K1837d];^SdXL1##Tf\
3W1cZ[GE=3P:_dL8OIH\9d7B54N]^V;DT]@0T?6V_^2JHEdWY+B-Y=Oc(;ESRH[1
BA5a<5:&HEAbD0AK]CA^HB?(c:4;E,GN;N>+3g:b66EHg9WAg]#Oad@)3X^a:gSf
SPc+a+G)]+KV3D<56PV7dP]=S,b(LKMC3TO[05?6b6/+>@S\>/>7c7d1XZ>VW,U=
+J:5(c]]PU,M-H+SQbbD=7XMQF(c4U_,]_B1G#//S,=FT3;<3D,2QJ#MI>(b_GO0
YJ&6#f=#PVXGcK;Q6&EN@d/F?f3(F3E0@.Zc8TCF7+L51-R7.:C@>A^6+COI;B7b
P=W8\:A87ZZ:(O<.FGU/1QI(2F(Bf&60C,Qa?J4aC[9:D=#P&La?YD\H>G:S;?.[
.;ZF]N[Z1,1^d_SG6#M[#8Ua.0a8PW=a);LDEI359?fU,L;YgIZ,bJ\+bXa)3#b1
d@a;6^=?aJP.^:+T^d[<H5#c\:,dA9NEYOa6ZV&^:=ecPU4],N;/;bM7<H?S6b7D
Y76KU74\?<^14Y[CU_6/[DbU)2:&RZY1gY4/PcbK92HS(.eKgF])=N@Q9(]@ZJAV
>d)EZ6HK\T;G<d^3]UU#);bR[,1EN&/fV7T5-SPKCHQSP(WCJg,Q^eM1:S@T^ca;
^T=C,g32HGRG-XL4F,=,f#(gTRT>#c6FG&FHI_L]A\A^gCK@0d?,^ABA(6K#[QD5
&2KHFT5GeEOB-\S#))GNS5c2>9K)3#>\?7\T_;c)]))[>8R/:?8V[GD;BMY5McG>
JXH7@U2Z,[LI/\XKD#:6D->J7U&N7c54Kcb9)(9[0?DaW+\\VE(KARCP7D<514\8
2(<C[f7P[[<@e[D/,IQRG4^:FC5ICI0=(I+&/]8C@0&[^CZ/RX5Q#gg<EXVV=PeP
[CeFNV.C8Q[)&P[S(2F]&7?,DD#8a5,]KG=Z6-eAUA\)JX1/FfOW/Mg@94\_:H;@
[A@28:-NI.0Wfd4AbP8(EQ/BN+T:GE?90;C_#gELG0O&F]?VZ\f#=#]UgZ2MTWMZ
c?X=;>#eGT[S42cV]#NgY(a/,--dYf2S;g#BQa@g9cZT=1?\1@^P?9#^GPYJ:R\7
._NX/4COU_?:b2dWMYT6>L9RR\90O_[7?C+&HD9?f).A09G3AU.e&VS-.;8ZbK#?
fPGcUOG<Ue]6MSK+4_gaMHT9Y_U>__8;;.80Z_PT7e?[KCKGCBG^DL;K#(UH2e_g
&\?Z-;&@30^.CMJ1;32KLNBefdFe8T)9f[)5TcX>.07=PTT0b:d^eaML]S[f24f3
H@(47,&IHeI?<@5\FN5VC<-D>Q#:Z2=d#YcW=C8+3eS_DP#2YZ_TIfO:#_L<NUVM
SH[[&_C3SBLR0@LLQ\eU#f<\,[:<HY16;-bH-3fBYNS=J6>EKbG^C1Q[D^M@b-<4
,([83KaOV\_V>5I<E#?=^J=S(bVNYL1aaZW-.WU3<8)D8.I]0Bd_8)TGV8HR^=F3
4HV;J6BL/8[GG34\I3T=Y6J)GG1(:E1^WL,U8=#VM_Y_#Pe1U;cQHd#Geb;:<6(f
[;OUH>c.5I7Rc(7L&b4g:aR246YBS1dAS2=.fbG-/35>S^b)1Pg,N:IDG18F(IFN
bLAPS/2aK5N<L[OHR1CV2C<fWP2eC1)RST)(E5;BY()D7=Z48eFXMeYP>9I13):^
UE1IWa_YBTF,VQKKabS1UGN-g:ZXYB4_C==^#B7/;JSE9)aR30^Ag=)#\MV5:PbS
ZH#QG3ZY&?</0a;/LaW=2^NF;^-bbXB5013SCcWe?Ba^EObad<&&O(56C]f68KW\
]B#3OK8@Ka\HJ1VV1I<^H/KG^\8X3>b7C:=a.de,La2(QIAS\0F2?DA;3f+EZ.K=
=&@]W,GC:g:,SKV.dGc-):+/Bga69B9W]GBa.^a79OCN@FY9c/g_#H?/\9,I46:.
cQ=c\:cWDK6:1E)9eLJ,Nb[)^dWL4>Lb?AfI)WEad?X2K\2FCYBa#\3^^F9K7&(Y
W?GO]_?e:(PB>ac7c95(O+QVe0OR+BZbAM[2dI:g]GRg-88&S@?V7.25@5P=N8Q2
Y7EWO1>]43)7SRg]^(4E>)LcdJ?.#M8JOU[=TR#5\U.R>X&(;:WQeY(#Y#AFO9W(
VaeZ^K\be5QOC?R=-C4\b0428b-43+#]L=LK\D3W)B+&8Og)WT?4K>3LND^CQa/.
=R)R0/G]A5=)?^OCG-a[#Q/RB0ZfU:DN;(_JeWLVR0@80J)TL#9HNVXY+9e?N^KS
4.>S:#A1HO6GEES9,ZO&I&&\L+KOI\:44adMI,g.K.DEB4+<8W+-VcD=C<7@JXag
G,M(GLaY1)2@&3baAU[XUfgEd2QS=(.VB=AddfVQVWHYCd5J>OQ&+fFSF4DL+gBa
#^UXBM3IA6@5Q&?0VU[44YV<MW,E(&B-<@fTSTJXK+58Ld@YBP5)&^4fE)ATX&G<
Mf;@90TUE_cGgWNX@;Cfc:5N=-=?D)G\QIeP(1fC<LFWe_?EQ&K5PaZO(WQWgdTK
+GW_.IY5),UEBd45N<fJB^WEX&0FTK@C?UG@LV2[_RCY(4W;aJ?J-FQ0:bA:fU(U
98X4dbRHTQgI3Q_g08RQaKJc4:Y6)gc?e85-Va\AEGZ=<3<:BLfY9-+^:-N26U^F
CP8-2#1L:5S6NB;YFa8?RZ:391Uc#S#YJc()Sf+HS[I7KgJ@4RFI<89;-ZE-Y=N?
G2Y2A+DS7[71BF7XWM4>DS0UQGRRE3-dG/5+Hg>2ATP:NF+LIg?,A7c+IbU:<@8K
EJ?K](bTV<3?_E;0-[12:dWG57MK3P=-b4^J4XT@[REUJ&C4H\+B1,M6BG#E^U0N
)<UV9#?EUU<->&L.a?g0K2\=CbREVS9#UH?)&P2+II-W\-Eb=M^&PbO;E3N>Z/DX
D5#L6[[C-gLb\JAALW4??#5PQcNb-bPH)Vf/G9FgL:6;5C=Ac/Y:C,dH+S<\+G#-
eKT5#NP8C5G(]107\ff8U\^P8ZS(+N/(YP&L0AT?a_B&3RUNW6B4fd<H)2QY(TW;
a\?A8d#JNBNM>F@V]ANbSU:)81eLg(O>\_.B\=NefP4IFeFQIT;a#Y.4IbOWY/YC
92DVCH&/?0MU21Y:AVW@TB>Fd_+X-O[MCY67.<4L_6d8T&4G_Bd=Xb>-Eg<KUWb+
+(VGWG#L3N^<Dd4]Y>I8__a6beISJ2MMaH+UUNAOGJM.\HR/,XKZ3=eM1YCN1P4C
.S6OEU?dA[F.():1V+E3#W=&)(E#(\+J97=FIaeRHJE_g\)4L.E@NC+#U)1a7M3L
#PWfNG_I147N+I=a#[Z0&45=^J/1_2/.f;bbd#;Q2#N3[@HEH)6a+-,83Xe,6XJF
@]Y-[GYNS()[Bb8^fLgg-X;E4^Z<T6g0UfUN_Adc#bO?I[NK+7I.b-D-PT+K]=9:
.F5>WBaE],N&;+Z2Ra@<=]#a@c?0R.)?fR/G]\4Mg3N)3G^R,<WF;3Ce+7Y\Ec)?
;Qe9(-+9Ne03SL\d7_TV7FU+5I4f^VH7RC._Me2,6dF:1>6_FD=D]f3&O3BaGX6@
?.1EQFga0SJ/S4QZ^72M?#V+IccSH;;:B]WX4gN3]a<IPd\WY#dZ,5@@c3JWXC[2
7GRI)8?9Q>Z44R&8SU?3Y?EMJSA&A&S9P)QK0;g4S\V/K/F7LI:S;Y)_cDd-(,W^
J5DgKSZc]](Bb)^0ZN2FFS(U5F62OUTeDFb\Qb9a):]QW&OYPS]bZCeH2:L=[Y)I
FcN<Y[69^RP(DL9a[_VM-4Y<37PPd#4+9G8#Ua+4HcJA+OUdS,dS\LJ8US>,(5?.
CHS29QcV4>F<]/P[;0BP0&cX?f[3]Q?P_K7@UV#SSU+36/^FJQ\<RCOeXb6E0F<O
14#A7<dD8H,J.VJL;;W[/N47QgSMEE9_.Bc>7aWfaE+)7^1dcB5V9]8T#5(Q,EKQ
;=M+>d[Q\I\Eg_B?S=#H<WcYZACf?WI&AGG^Pd/\E^B\Kf-&Q2S7?afPL;LI5gM\
^=#3dVP/,VYCGf<Z-ZX3BgCGOLKD+:^dC7cF?/BA>KF&,9TB0dF6_F#;X9IgfbKY
gVBG;;6cRV6L-BHI[&\1N1+31LQH0M-5P(d);@gJP#W?8&6>.N_Tb3399d\QgcZT
2bfbRJ]1GSdG(P7@TaLHU5]JX]=73+K7b@L4P(-L0OBaYced=fD/LMOSOf<29U/1
.bV.W?SF&;U:7(=U<U?AM=RYC4WbNeK@)N;A_S;/B=-WNBY4G__H-_)3H6UW6Z.(
2Q\A+f)&c5[&Jc(2RA1E-2Qde3RNPN^=#X>=96M>8M<Z\^A7H:&RFL_AbUD4,(SH
O#NW(<L]f2e@&=^ag\&ATF13LV]566WgE&GL\:),=6W=8&I5P5144f<<Bd1W]cg(
R(A93V5cJ-50_e)E/&/_3&[5V5]&:?YY2I6@D.P9>9F\-b6SJ2-XeW]aTRV[2d5I
gWI54JCSOae#&X;DcVM[d&)a+J_&-).I6P/WAAfd,Ab[N>>f6-\5P393f)Pb9KSK
#GJZ)LSR70A)<0]ec)gH&B5J_7NG1:ag,G+F@P/ZYOQNNP+1:O5__/>/c7Q>X:GK
\^E<C3WUBI7A^3:<DAFAEMP<5QU>_d>7cB/MT).P\[>TJ_?SJQ:&7T,1;KHZEE+F
Gc:-W8LB/8PGL&+2.41,(1OgdGdG_7GUg@HY\W;5GBW#K][N]AYR69RJDe,>JH_L
[Af?=a5:c+>f[F(LcO5dQ7e#>/#FPc:b<0@,8JUKL,;,81MC?>[e@bRbWLgABS6f
J2&I:KPF5NXW8V_T\;aNQOMcDLf\D[\^RX0K]5UfI0FGW9D>G=+2O?O&a-_CO\bA
YJPW)?JHF7Y\^Ke7X\-)>;DA(U2_FW((7)+EePO)1U(TJb=^Kd<)GFFIR)N^OU<A
+b>7/_#GT16bg2R@&K<(OG[.OLG]N(J:YC1SLegaD&86@POD2U.&Sd^I(Y3E93?X
CB+93gDNZ,KZ]ECJGb)M;Od8.P:C,4B>SVM#VRJ77/Z);.b5UNVIWVE51T5R)c_)
F;dH:45O<F<cZ8BT(OSJ\4E0Qc1#GgZ7QDXGU^RRAZ=AMER]4,_1KKFSZTO?&2Td
.0Z;PT8DecHd?aRPDH+7edFP1Y7Dg[O>E/<6O^[OO(4#+HRXfZ/?SK=06I1JM@>b
5PX-9?4H:DW<a)^cU2Og+IML)L>9<]OfI(9fPbDd7R.8=BU]8]eU]gX)A\c7?R<?
Tf\H)W)OfFQ#[[-7H:G=g,LXbD)bWe_K8J,&9Xg6)45R6#>:-D6^,5SdY\0)&fS+
V&B[M1GP(LH81f[:#3.YW_>PE9MS)/P,e;2f;_V,NP]<2g#+]<Pa]O^S<Obd_5S\
b5Y^GPFFd,)H9=43?/A0cG9P5W4+9A/)5MO=H]+6C/-602=PAM\5<U]1OYWMe][G
AUKP45Oee9HS8L@ZR68I3N3X4M1Lg0.g4Q\EfT<GT@\Q]NHbA6]&R\2F<;PY5;AR
?Z7#O4+LNXMGZ[TE^I+^0_KQe7)]-Sf&A)N/EeA=aU32JWO&f_QefK7DEYQ+X_:^
]La1J[,VGf:P8gE\AUG,J&?XRO64^8=W1eUZB8NdWFa8\Y8C7@ZM8OI_MK9V+U5+
PcYVLHcXOaPTI9D^37:R-39Y;/#6RU4ALH>JUbRZ[7bQ49_3N;Cg^Cd8\@+.F4PT
&S5f+4bNP8QE@B3g1I3PaQ<9^_/_52G;La@4Y3Wb,PT59)N4RFEH_HSaC4/7fS<I
8Y<gdf@HAG]B.#f)EVHH7JJ/))G:4,[AHT;LU=e3IX2d9A@ACQD,\0ZR)3J@AJ9A
Ib_;@ZH#&aC4fc+Y_T1OWAc>&LW)bQRPR:W=1DV-T.(2TV>M=bFO_A>F6P7#^Z3Y
gaB[VK4>4VT&@;Hf]UNZgaE=;I]UYWN?=</F#;/_+9WHP/)&9>bc@C=?gCW;1K4.
(T1UD);++.\e6IK2fXD@V0.0^550df)+RV)7b6#cKbD,]X(c)KQ6;@MRA1)WMEZ1
+I9;gTFP>Z3B,_PEZa2_:]?](O?5]>_<:M3ST[>g0N6)\+QB]6g?1ZL@g:F5L9Lf
1\a)EGTOdQOAJB7-geUGDgOg3N)@U11_]8Gbb??@KaF7+>GJeC=64D/AF=NDF6B8
[)LC/(^X.(:2N<1bYUW-Ya\gG22X4I4;+g89ZTVCe?9Y0V;Q]^6Xf0bTY:UE69#M
@?=I+9L:.[]e)&dMX&O7Qcca@?Z[FW(+WMS_d3GT,-(<NM50;<CL?-0;f1)8HHD^
)a@@X]g9LN5\)@ef0bXZ^@TQ^F8E)/<6+I3@Q1:P?EcS&_DW&2\HLSOJB.L5&-J^
L-=):#HG-_a\W0a1e#4R#e.TLM(>9]H_-VYJ[>dOfG@Z1:#)4/ffQ]f.+XF_a6Gf
CY>EY>d17=LbF6^/]8-EV=1TGS:V46D4:DG8(cKTA/LY71dcOb_A\]5;-=6F<>\B
2bYF+_]NfO>M;3:2Q=967&7EQ3_\56d@GOWd<E^51IY3W0OPWV:gB7&9UM:QKA41
NO+ebC8&,BVR&^6[/\8@)BH_a.7b)PF>?2)T4B=Q@7CZ2N)e+\M1O.f8?-OCS:/]
H,4A8<KE=UbT(OC;<H.;X]\BF+Nfb4#Z9;,UeNS@7DIP-6LN2A8cCagb2@<03_b1
?=b_gS7IRc#V2#)?ebD@MP=/XN-C#3,KQ&&^7KcBXI^?VebE:Gd[/1;H>eIXJZO]
eT#88gbX;O^6I9a+Ia<1U7QQEUaVQ>Ng^MLC-#[\L86=IAE.Y6T&::?8J-7R/TQE
aC+gfJ02b.2c@<9g1:]cRE_5B(J@,:ASERL/OT8EHQ<VT=+2&PHM7ZP^>);O]#^M
U;-OS1\DV)1MbgS?;A6PgZMY1=\R/-bE)cV#FK<[d)eE=B4>E;8b.85JeZ@d\H9d
f0-#,9)bDWH8/f5LK.,^;=[.XYBMJ[cSL?dgdHDJRI2f56]7C--cUKVC^>4V.C+]
a+f;Q[acO:>\1(&=c.TB>?,6DEOX5O4,E^DK&RCCH9LZ^A9e:^Tea[=YUP/+:g,>
d8AZd,W,;9N6H9KL1Wf^C,SS)+)VUYd^DQ^2Xc?E;IUKRCUSIOU[5Q34Rc3PZBV9
^#)Hf?+f,;b0C^^DD,L)^].K@TdTRIV>+(;/bR?K<9M)^GWE?OSOX&I08O6Neb5b
<(?U5F^a_@&R^.HGcJdXOR0S1X>Z=c0DT]<bdD5E<TMF4dR&5V1E5=45]^T2SFU6
+ZP9K06GccDIgWXfI7778/HFX#^>1(UWQEA\6X8ZAHR@.Q1E+LWFEZX54GgfD=Kd
\&R@6^_1\H\eER.357T#GI&Mf#5V]:?+-EEVfW?,[2d.0#9cM,\>\GDF^]A/6]\E
L+Xd>cW8afO)eV51bZ9+abKO;gN=7<_/&Vg\fU3DBDD]]JQ[Q7&>D=I@MV8,aBd_
dSX4GBI(Q-c^U-0?cJ5gQWSTI,?354afA[b(NV#O;-&<6.7W6N&NQ&--2PA3+5KB
]Wb5>?D3_eY5L]TUQedFCaUE5ERN]K]K..2>G\^aSMV,]0f^ZKdV3=N5E/6V9BBC
)O@R_d?M;[_QWY]@#ZfZ;FbFUa_VIRU7K8P0V<?[ZcQ#F.cYa\&]<eHKZ)S-E:D,
9#55JG1=AMFR8XW]-(G7SRQM81+.@YK?,HcPd?S,/)D/L=.O9Af^Yeb4_/88g];T
[5bdJKRc>_.aT++3;SC<C6O6;GX&KdHS5D]U2@@?ISDfB:<aN0A4e_]HBfA4FSLP
K=:U@F[dTY=GPa>=X_5TB>cCFc)f6eea12X,PeVJ1?@7&(U:FcF5gDPQ^J?H>NAc
Wa(&EP1(+L3,;f>VcA(PMT#A__<JQ>5P=C6FL1>_aV2+X</b6J:K)ADSXM+KX;ML
Z\W9>IKL8cNb5G@F:cFF>3db,GU9F?_>g=O?F&6<9T4OI0UD]V2?JH/=7T;cg86B
&@OcMd<2cd1I#5[B3+a<=bKT8F7QFNP:ERf+_LT7e/B&-OW?,LUHe#957J2R25Fe
+YO&)>?TRG8/U<4B1[/VXa:A()A?#;5[)=4?D&C^+8@6&+T9P][?/3(-g+1/VJ9b
0Q_U1@?CQG/<6.IENBEA7UGe3=?a^?65L+@==NO\4GZ8IQ\QHbH:6a.SJ4d7LJfH
[g;-U^VZ=6/)I):g0[4F[O0FQGg^C[<_NBdc&;YeX)]CM(@7EFO-Q;QXEL+3^)[E
4/314LYfWML2I2S[g8=cFQU+&SK(XB[R#E&TRfC&0GX.>3CQZfR1;GH1(VAbOWCF
/JD]>8g6bT;VgfH_]ZV</6<A@H6/F,.FZL:C,dPa\H?f<b#aP1@DJG[eZ;DFW_Be
Q\Ud4PV^bb;\HSaQ73eA_VdE(<b/FOLa-P?^9PY6P>-YLQM?]8aAQJTCCYE;9M?F
1,L#AY]d25IW/);WTXE/,N=gWJ^d+.\AGI./&^0-:4O;>?d_\Jc7XC\gA2\F6/@5
J][I83C6cH\WQ[V(X9?>NTN^]OIK.PY0G>E-?(VgXOG?O>#0#[S?+FHS>B1H<R05
ZNNQ4/PCBF;D<T.FZB&gTIR,H+PJ[HBX8O^A>PZ6;#Y)F3.O>ce-<?Bbd:Q&)<X_
WEMIL,O;a:P\RIED1W[f0[a5RO3Td+gN1:D0;dY44/E2[T0a1?OZ;)S5aWDH>I4I
KQS>bG?f(a=FAS.d1<MD[TK=f2ee68Y.AUfTKV.f)YP2HE>c65&06B9]CcOR,_-_
YVAcb=,;U<=e?#G(H?^?I\@JcJDaeW+LZOI@T(PZJ[8aTKZEZ9/YgM^^cH</I0(O
+7O3O#+J7HfLgIS295X^]R0S#EH\a92WYI(]KAT]G]T4E@@=1<?6_@Be[?I8KS8I
I1TTY_>W7ZI4Y\.WP(da;]bR#SW5<N>H0O4&CJ>3?#&@^9A,:#Ec1T;JA1HTM^)H
X2FQHdI5RK>d^OH0[,<E?a?_(>M=1-]E5W_4._E@Y=O?TGV6(5;:ge59]9U+F(W8
>Hd?<.YK@:-+2T#ZJ?5\>4N,RfEE<81-O,b5e4A0a-J8&d43\_<e#/>WK0[Uc0?X
&RaO><E0YH([1[4:;cW<0JVf5X,9dW\V&[(5MQNIY1V+I?M.?4@96F;cRdbAbU-a
QfO6-g2>3H>+aZ9CC-.NDA+J9]]MUF+DcWE1_8-I4M_TdL,=W0aPNXL6D:dSDM_E
0>UZ->IK0IQ-OAAC_#7<7,M9g.S=>:I4^([EY\^?)-^9X0DY.<gJ<#K<gW^N5(MS
AL33G6Jf@:QbI.5YS]cee2D.^+T:CFN\bHCM9E7RHZeR^a4b[H)CZPXYE]6b1Ua\
A+&\T3T/JX)J4IGK&7C@N)B<(XD6:D:.=<2AYH05+c1_S,4I+,Q?d?Q\;G3B=&Ie
FQ\]MWO.EBc37L5EXQ8#1W54,We@__MP=55Gd+:#J5U--<I23;DQB&TP7&22HX16
D3LJ0Q=bG(g^[H:@Q]e43;YC\aJfRdZX&<e.HCIS_W.(0J[df#]ffV:M7VRGe@d)
fUB6?A>S1;dW7T;]U53;&[P],R]]NSK2W<-&9bCE)4:fLN^KZ&MRT)e6OIH4^C=U
5ERJ&=6C8V<&TGVYf2>1aN,.eYPgSAWA(NFd(<9@4H>^;UBF=(Y7?4I13Xf4O:aA
J0KR<&^@IdQ6M)aQ:2JLCdHGC/G-\A__Q>M+cg7TdHA&I@W0<V=@[EWFe_aY+O]1
#8UM:2G)L5Tb;^GM6H_92TNeQM@RC?HE++)=6;33T@9O\87QMcb=+:TAFFI43^\K
6HJA;7[W8IS:/6Fc+/]J.P_^c93b5^PcN9-J6N9N+J^+V(Mfc,M#I29M:XHQ_><6
?.ETeEZHH@/d\^O\-N;gc=;Q?FbYag-F>E#[a^:Z)&MKfG3FfbI>_Fb5#Z2GFb=&
#1IR3U[A0A/.fDGT.=.EegKH&MR8M6U<96[f3b@Q2f>,c8^FWE_I?aTeaYSWe)(C
>MVMG87cUMR^>EcO=FKR(==1IT@(Q_HB#5f4c4/?GF)^:,=G9+[I>a_8N5-.V\R?
HF94]@=^fNCAKGVHK[3.FTgGb\2c=U@9,#-d-=_Lc)PZUQA_aX2W),Ve7AUB31=a
1YU]W>SHG<9S\F=_][G\[+A=@K+^IZ+.&7PH6JKb&a\VL-A<<A3g&\/Ga7T>UWRS
4b(/RaFZA\O8b[?a9U&LA]93#0W>c\L[MTU2WSK0OBNW=PODfEJ;-@1_Xae\C-If
gM=L&\V>^=-YQ4O-4a]GRMF24_6\aYN987\Oe;I4O;[.W&>H+834L_OGQ[EV3XE>
/>V#C.<+0eY9MEG9N59E:E89TAL<A;84X>J\W>dV8I+gP=:[(_S[09eU[3PVXMC7
=?QQMTRH4K>Rf6CO^[43?Z4_Z#bE40_=SZ^YVY;_U02TY83I6J2-RgD_b^X_I.@:
H;>I=GB(O8#<4=_A12R26#R,LQ,TUYS.0;YIK=OQc)ZdeF1fN?&</,f?#?)SV[?E
L+Y.E&-U\bY+/:[a8SAENRe8FHO=B@&@0;V)Zad#7L6gX-+;-g]&2LHP=\a_gfcf
:H#O)XB:g)1\MKDITTS(107PP&#?e&2_>QW5_UbOgeCFWSLHS\1X.R[T)9_LWdW8
>VR>]),XDXf4X/OK-a[7fQ2(CPa/DHfB.RR#G-3IEQFaMW1CD8\2(X^fVD>O.(Ud
0QS1IFeMcU81M@05>KF7P)/QV>Td2?)D6<-QfO:YM)-,21bV(T3)@26J779]c+KM
A/Ua/3?:V.Ec]Wc<E[HI@8ZGe.Y3NG7NEK55)LY0YW0>[:e0S)H=K]](I,#&8?Z0
CQ4K60E>EBHf8dg^gYc-0#<&:+BY7[]H7;eWJYBS8VA<S)=-N]0RBJ,HcJTO>5eK
=NVXKX0?e3-L8d48&]SQVB3Qa#.OC7FL:Q^Qe^\;I]]]a=7]O2g:;S)\L0.R:G&\
@d:SI;Nd7E4#MAVJ9T92VV+NC/W_e1850D<e_J7_fSJa@./[ZNf)DYH(\ZUNOXJX
G<B6EVM@@]f>^9M8XMU_KABC<dH,((-#XNV;TLaB#4#O;7a&YSb,4Y2(K;Ya=ce\
B3[cTBCETWEQIV4HRbDX+;/Z?f(&-c/FQKT,HJIWZHS-aOA?fUXa20U8I7=a;(1J
4Eb,d-e>J<.VX1XIXDSW&Wc(IC.ZJ7TZ6QWWRGeI@:.e/YODC&EI(I:f-HbO#bL7
0->2&FSV>bb2Hf.6_-P-9@)(>ZA_5Rba7TY41[+ZV,E&4KHQ4f]SPL#C<TWQ:.SB
bU6b6/ZK_dVA]NcgTO;3S+?8879JL@4&GBdb8#?gbZZcJ+A)0Ae;A2_&5VH5_+Gf
R>VBW4J6C4+7(=B+Qb<Cf6BF/&L[ZT73)5c963682DaTWJ)G92@)c,9B.KSPYEe?
d\^J@B.;]#3AIa14R5g]L9:RS1LE1cN=/AEEU;feA(0a)0KZ+SC_Xg(gXA+)<&GE
?.77S61Y(EQQUOG,=CT_2a8S/[5fDOZ<>C<7g@F,47<W,MU(GA^1<\(WEOOH(8]+
YM]5JaPXCPV(fV-aOa9#FKVH,3@05Z@;=1d@/,V8Wd&8&M@689\c;T&L:I#\cBDR
dg);=aKN;UJQgf>A.e5R9BJD<4<;TBL,8dBQAEZ:5#?\8ALST[I\2c;b79M>D+L_
N.Q@CTT#d5]BD][LMDZfKX#JE:\ccg>f:QKE+<#f)1TYZY&^e+9-cI1^^GU,JQb1
(\?AS#<8eHGF99/F1RTIY2/G-#7=VWO0P]#S[&0FCQd\2b?>\;\A2;H4_9;A,c:N
<4J&Q9PB)^HaU]7D,,A#b(BAP(=1O2YORCMXNXC6YH\G^74JfEAcZ;-X.bV81,VJ
M@,[CV@-S=,f@Fb#^+2D:cPeHeXF78QSGN&8a1VX1V;4=[[Kc:>>[G5V;P06Ja\E
VJID^_GEGHS3>5#aEH:EX(a+f\#;#Hc=)1-PI26bVc&#EPQ<[R6TV-B3+M@0-Q7,
R(eX\8PddY;-1LU<-7]^,N]=0f:=S\VS;J(6#b9ZP#bP)H)+#R&,F=Dg<b;0Z,Ea
^cCQ3C[&^3GT)@Paa&)9M3P]UeU/XS;.->F7AY,/#8/f3[&__QHMb)7<(E6Egd6]
H1SdT6SE(1HaBKeE>AV-(9U#fg,GS:WBbb-:@PP-DQRN_]A^-U24)-Z:7;(ZS.65
bG)a)DX:g_F-S0K#dc.#_].A.K-eBB7e(Y&\3bST#Z>0dJ50gZN[6-\6<+UUb_=.
(MX][Ae&984NM>POZSZ,cEW.VRHUW88K,dA7N?<&^)^e]gF&/W\;EC,FRXVbXK,A
?D;a-D]R,/)6-L;dND\#Rb4I89?fH2YXQC<THVMN9L;GDDC,P.BU5d)9.=:3fTS3
1?C2]&UOH5)H<#^;5cV(LRFG.5WD,<0Z-50Ud2(6GDCcS5I7KT)TD:RXW_IEQ_(>
09>^Bc_G[ee9V_:RESNf_E?1a-)AUIY7PO1eJ-9f9TNCg9J@;PZ^ZWdB\U<X5<da
)->:f@(>R;H9N3;^^0<44Ne<X^=cMP?LEXcW3/8+V32RU-F5E7dF589Cb_cZ-LX9
[Ucg//WF5ACM4&A;JN;@W-K?,b@.+^TX7SBEc659;bJG<4b?[<QV(UPI);KE/:>#
/6,X7C/F=dSP78:^=_&4W]dBbO<EcZf?:/^O<]<-5:(X8I=VWSD851ab?0\4Ab8V
308bL3_OG9LH#?Q:O?_,Ff\?6[V6I::J>]UYT]Y[@_3)1/-HGD&^d;[ZW^;XK8KA
##I-N:1&_O44.gQ:1;603RA.P3)1ZDTd=TKV_50c9JPLBe=6[+a+.:C.4,K4^&@7
CXG;^T[;9>9//?10]9K]C..gRf:B3_?G-.CFUaLa#F//,;8gc2aHITNRfSY8W\eB
e,]#NQA+gJ8QDW)?E[V-<T-M<OM+]W,(2VKf^3PW7DOD4_#MWbNb9\P;EZXNf:#R
TYc:ILeg3Pf[3]34]W04NRTQ7>J#=-\LfffgS([dYYe0&ASDDZOeKVX8]KF;GX.Y
D]V.)Y[G2(SeM:I5d7?9Sd[KQ89_IDA>(<abeRFG35c8[VbJ(V9X1XfR/GUP-cJR
?SB]0RK+OSRI6UMb\TB1XI0#>cG2[]OTA[6-5<D&C;]G=ZQWc6QZ;57P.QFAB6-\
@Y3]TSd.#PE&+A)VgPBQ7U:6DHf)L3=dNCX;&XWJ)T:+gKP;>WZM^??],LSRe[8f
WDQ?Q#4Wb>^1W0GN.Z#Z.O\O\=Vae4C\e_U2aBfe=7bIGA@,A0H+FQB@IEgCZGZa
a0O#;8PBcHGBC.0\+\e7d6Hb\/WZXA1+E,#YOVNO/PO=#H[?7EUeR-gXAP\cL1[@
?2YT.NP<9U=:@&f.N/;IZ.a5]SHJJSB#VaHfOPA_X,D8,V8.@(X2.AF,FIdY8B;D
+bY0=,3fgcJ^5RQ(N/./Kg@N7+7J>S^/dBc6gcPCIS><N//4^CTVVWF&;e]-;;0C
Ub5dA0f<ERM?#A=DBWVP38a9<L2Ib@,0=Fc>:9?7B]2bBE>c#d/gc4?Q6?E5[VgT
J.JVQVYO#fE2Y#O]HTSS?G@;U:eg\:.<>bF9;Y=-b(SO[F3NT5&_4VZ:+#O<9)1d
VV3=M6Q,<,_EZX(_3+64J]O>>8OJR/2g8TTH#8FF>Y>]KXIQd#F\UQBW/e(NaPg+
>?/D/V><(ZHBBO(YOb>8+_KMC]20X8OfQ(\9G>]G1LaII4DdSL^;.f]c[8H<VBLD
-<d>?H+?F2WCC+L.Ygc(TL8HJ81O:?\5bN@Y4BQ6:YKFa:LHB?a[VZE8]R;gJfe&
K\]Td6e7Q/6C=GVCND<b#<1_HY9W7XO)]IG_\:Va[//>#WJcV9M(@&fG4fIRDR#P
bdY+;G0T+eZL#MKEaEF\=]5gfOAM:Wd&(O,Da72>L8Me@YQ51EXVDXDM8D\D>e\;
VG+;&CUfZ61TZQ[4JR2TSB[7&DcZBNcKL2)H>]NF^TgX?-FR[Q/IW;@@W5SR^X17
NOO3,1edS1Rd-PWAHA87a_5:8eG749(+NC(-8?L(]DNg0KHeU;[VW@EU;K@]\=)]
\NH?I2W=-E)@3;]T?;_:&G:I-0Ac(Q[bFZ2<)X[3+])ZD=DdPb^574^AP--1,?J+
)K0(S_249BeSc80b>0<Ad0M<9Ge-?dVb&8B^&OZ5XgOJg4cHWIb&a9dR0N=&6L-1
T-<(,=@Mf4@RPX=;BP3<E5\HU8,a,U4ITVIN9dFN_c#AHQOC48/=^_G]ETd1O>LI
]^E(,YES7:.XZ^L2d^X_P=5PR]d]Y>S<:]1\&V;4b4#g/W-<?e&R-[\#f#U;LeTM
LEP[Y8@(eRCee(G[>YcB](4S4KaPB^e^=_U(=?)f=U.^P(bFN]&UO:73X/ZQ2AU5
Wf;daMJ>SL<b[&VbTd@4^U#TEAA;^@-5B,E@C18.@Gd>>ZP798g8[VNF6F4,1:Z)
UMA6Ke/?C689IA]bFPd2#1D/0F-;W8UK_afJKL)NE4GD@Y_=6dF):_&K-.F\I<aN
7.MTTg.MBDg]?V88T,4I?1Y<gD9a&(W-7-OS2]1HeaT6>/->PG/F<:@\3Z7[IJ@7
A.-GgB_d^AHSRDZVAH<TSXg<]SOL)#AOA)B+e)^b@N\\?^3A&cL=Q<UFY)(bF2FG
1?49H882Z_GaBHec&:.eFXc)/@<4M[72T0/,55Z>Ie165Z;P&QNPaQG]e=TWSIYe
@MPg)F)<1XPd,9JXMLc1Q5I94BgS^I<;Q(P^B8SNP1^cd5W:\bB1R8R:,&3VRZ,5
fT9CY>C#OG,)Xcg]\2g9<<HJfN)FJ]3&3=#UBIT71@Eb\RUQ/P(9W,KMW8K]R)eU
15Lg-+)3&GMKQ&Nbe93:1AMM31?[:40?X-EKWOQ/M4T;O/dQ>TG3,0Q]C[9U#-Gg
g8@\/V2U2ZB>YKZ(@GLDI:@Nc?8#)W)6c9@;Q_0U2:eT?MQ<&P09LD2gT8W?3HAZ
)QR;/g]+@2fb^bO:OgEGP;IKT-3fXMg3_ZXR+AL#.J1+)c084;@N]P8ba5GdOJA8
C)<g-/b[5+I3H4\#fA=ZZ7#>[]D#f<)AL](,O?4((0@V\B^N:aU7BO]CcZKQG192
O(J2ZZ03Ra&dUXJ9U6Cg5b&/RK-V6Y.6Z:7IP8,Y^-UQ_&6a:HS2CWC7<J6\9:Y-
K0f8J.#0:S;4D:(,Y[H2KXA<QF^T=Q;T.2BPb^b\UAGb&,J3aIE?>,;f@BM><D=A
U-N@=e<YT]cP#8T+,8B0Y>WN+:bEEJ5=PMcRZ0Y,AT9#g3HK_8MKReC9]SN/,0_O
SAU]JH<V:P/L><:2IQ:&I0bD[HMEfg<#+f1+/EEJ&Gf0W\02\\3gFC:7N#?LD/J#
B16^;gfa\[Pg1V;)S@V8\bD2d5,a?MBcFI<?d-(X6a9U?&#=6;VRNaGPfO@9U5<=
3QbJH9E+\TSHXVd9&;UL<1X&ILSNVEH);3217-O3PW,7.<V:]IGO(XO+TEYYOPf@
Eg;W1UQcSXe(ceN=@FHMJa^eGH?RP2:V>9=9d@34(cJM=N4=J&;_2;BE#HKKQ4=,
,L&T..6\QeW<T<F@I/:U=3.B(T8SI1a#,TN_E,AI3WF(+\P_URgOL]=X_,,U)7@a
]O5QU?9[VE3EQPV.:Hb5W:Gb4c-Ccg#0K^B-QIXQO2Y6]-[WI7<ANG5&5ZXW1D-/
-7UIace#QX5\dZHC2ZNP@_6+Ffb_3(,F:-/O\>Q-#)Y1YG[<(9Y\eB3L\6;1aJ-R
_E]W#V#JVT&?6LYYPMIfI;XUe8-J/:V(1\^84?0O8Ad5A:WfP+,EN,Z==7bMf[>=
\NO.HKM[^CPM:^KFZe3X,bfLgSH9CK96<XPHcU3Db5O.5FeW/Q;be.?5<D2CFSdf
SQaBTOKd@9Kf^]RU?6W5HCE6a):gO\,C+Z+\5K_(EDLVQ,IV&HS-AAL5KKUOPc@J
\/[<#5FVY:]bHF\,<c#De+KTg/1C^6Y,D?SS,SB.5d@^#cM047WgSL/dF4OLWQV?
H#3WJU=Y_?Z02-^=WfSZP.]dCBb)1_.8E)HZ=+=>V+OBSe4fBY:N<\+O9#6Ad4DC
9Z#@GTH)XgB+DON@L2Jc_J74QDDPW>M3B/9K@M2Z-EX\V0<QU@#_QP7XJ[&Mc^&J
M@)456K-X@RRXfP2RKG_Z+<?W/J.;BEYd7Vb&Y?UCNM=KRK9Fg<LL)I=.eNT7L)I
XBAZ<LUS[-g+f190VS#EL[-0Z7RZU57aZ>H:);>LLd];/\07&R2KM:IF.BVL)O&c
6>b(U5U8b.VN=LZHK/Ve?f\47C\=U.73SLW?F1:J;fA3#VVFL4cP1^221__\JQ9?
2T\]/:_6c?UH@VH0d4P1F_c:<)H;_9(R(712KN.P#SS;L_.=HcNf(fSb48Rg6[)1
7bMQB+,@VRTKQ4T;PC2HZ-2E?TgGK1a3^/MGIQ5I#Q/E/1e?\JXT[#[65E<<[-<_
cCRY?I)H^XIE,I/BU2(+L@F^9IIWT2J86b/_W)?66=g2UM&4MGIWI_^5\cFCPB6T
VYE4W6->>AN6V[_[_49ZOaU_bf<X9QJG\</Ha(.Q(;GAN/X\PdWR15;2K?M1U##R
CY:c_+M6RXXbY[C(1W\)A-gZW6;_?H5A.91C4b2)UULa2SY4U+4)(I2F1F.H>YG/
XL0_-J/@0eLWWeI&GE7B=8AcY)3NPXSJO\8;<e2fBD;.L0ENE(8JNJ@eg\.BO:3X
EdY.)8^+aJfEFRO94@\#Y_V#TDg?2a/;NUA-Z5Y2)E[+V0\I&8DG<-O;HB^1,(bQ
^OY,g>1Ge\63.2(1CA6T<6-^QcH]P<:T56YbfJ:].EAY40B.PDB,b9SKOQ0:[)R5
N3[(+&Rf&&T017>Lc>R(SSCVP2X+,:[-gRZ?<Wg^2M7PFUGf,5fWaDV\ECc50ReA
Sc6eL]D03A1[_C>5<#WGJV.3IbW:TY6=Q@)6&XBQ.&eO^)_CU]@3=4_-9M#;-.\K
KS^1+:cE?I2gd_4bE9;KU<U>:^]NKCWa8UR@+.Re6d=?;aEM\/>0A_F1M&a78QTM
NE#^Fe<GL3b/RRabI]QZN?]:+X08.L7-C;3O[Nbbc6_-,<Z3R8(><,<F4@<K3+]W
L<\d7_U(<6UBUZ=B1L;;@)?\RPW)9@5CJ@O?[4_><a#RL,K:.#/8-S\9I&O3.V4P
U0)CF5?FQ1WCZJ-fOSEQYbO5[NDaG&P):U7SN[<)CNB7S5@=^_b>8N7^\W1=7<gG
VQ.76;NZQ4B(>M7;Y)I1gDJc5TfOIgU_[0OZ8+ZB-_?2cfW?PTf_2QX)FD;D2K&_
[+=(76ILQP&_YZ1@A]@4UBBA5Z_8RG.UQX>Z16;Qe_:=a;Z@F,C<(aQa6\L8\AQP
X=3DLQ^.BNN>:UR_QZ]c7Ha@42\&35YNNE]cdU^e)O;RB[.(&T6^Sb@>d27T:-1]
+ZZ:UAEg\g=1Q-E-O\MbT_fCUU__L+IY.ND4d36#,)bbE9VI\.EUEN=geV0Z:d\9
g)S1H4T,3cHJAe>Q3f?^E\3Fd@R_S3J\+M\ESKZcB<b9@Lc[2]M2@F;[V.UTPFG@
@_b4#T7SQ;3,9XNGaT6f)9QEN2,=bK9dYQHfQH12?8K7<^Y=B.LC\+3&UHa-OAMd
0=D6WC=O[#U]GRDVS&McPRH#6V\O]U(bG0HC)OTQ>RJXE>,G:O9S1_X[(BM]+dVd
7X=8J@>ND,MNLTUf(Yd6,T7g_9>YM_JU^4Q.@<-V08E>M?UYQZV\e-<Ze-e95I)J
F\0=?BJQGJ0g&X]\aC++]5P6f:.g)CCGD\:fbM<\1-<6Be,N\XNPN/@Ac?5fZMJ<
Ad2SHJ,VBK^BJHMPCc_@f^YDTcM]JW^2fXfA5Z;,0)=b?LP0N4PX;YT;62DWgbDK
&:0\+,QN2FFc9,H][2@5FZGY[3Z\f4;+(K3g9T^P<2PRXJGNK[40@2bb6N6/Pc?<
Rd[65e3/NX,>bC8fT)(bb@M/ZW__XdKU;F-O^?,FR<B6-30c_A_b_F_\H7\BSWR;
-f?fY?.SY5M,?^XBBF74F?.M(g_#LG1Lg1#B6fd?<,1LXcgA.g-d,>NF33d);F\f
b\M-]Q6NHK]5Zg[Ug_=,XQ97UcL3d07:1&IYcE5+?V&<OT&GJ>e]78\SE;&1Wf-(
M:0E]55::-Y)/>=SMI_OK)QSF&^H7^OKf>,4LW1UKO8+@dg_1R2be:c)PF9b\-8E
KYYc.@WL;)eY&QX-<JJ@8(-,?V_=R[CL:]6G85VRDJ.>C_\&\ZNK^e_4)<,AQDO;
V8-(OSXEWdX[6^,f(RZ(PLWOcWD?g-PD5gJ9_VFbbN3eGRQMT?CYZ)a=&FYJ5V.:
b(##\1)ZDT)_TTL3P&2DOBYKF5X=Yb?J.&HWY4D)Q=7dOb=O6I=M2BPTO37g-E9#
AD8]6>X;?#:#G\9^8CYGPd9Ga\L8^U7Q]KVG<?eV\NL/L2G[^C6Ufb>+8\RE+ZdE
<Q/^F]-CR&L396AE5GGFfc3Y\Q7BUa@/_NeOS]:HDf,R(\-;Z)9VE(^bJ1@3=H+<
4Kb3)=fE378.T(?^7<24\T0cV)G<7>)[XTI?^H93J@LFDF98Q]YFT_+AeF]3fXdc
&_^KW4GCUV9dA<N[(9)3Z;0P74Oa1P3DOB3<WTK5DE#=-2PSE+IZL/R?-D,<O[LJ
GI1K]JRPX7eaOSEf>0+X7GfI]<.<L:(_NS\^9MEL)f9WV7#KO?b35La1E;+[]=X,
D;S?75Jc>RT6KB_IU8N-1O<6<XC8&fI]ZNC35Y(AANcWEd7ZISHU7g2<=-:Qb1/)
+R9UIBHD^VB7O[,R,)9HS](c>73SUDgK23</=52[:+ZP(_4,AW:XbRM4KKJ9?6];
DSSY]F7b:K8bb3A,UgeKfRP\Td=]7Z);-?VM_])6S\CA4Zb&68K[I838IY@?V]^I
)c)X1;02McUbHICI+O>)2e<9\]_O4FK[[6:L;;,XW9bF4?ZB&..=XYEPIDG,J2cb
d8;V2a,..2PC?;aQYE-CADY,@=,g^3#4:A\\J15L<K&)A:(^^d>b1EfWKVe:&?CV
>>>K18:ZVG2(Q)T;N&R/Q)0VSKJ=+[XH-.f7I-589^>8:/b@FSVD-Y=?>b.?BWB<
56L:8^60Qe;b+/O<6GZ:bd1C-U=--N_dGCdZ^-aaaSGQ:fQTRY\<F^?X+]X&<T0G
_3SUBf4(Pg^QMg,N2Lac=<K>XVQG^P2^GI2(H)+^3g^Of0JEW_NSZTbUI0O(1c#2
]1a_)1FEBJ,U-gfEC90I:Sg.gf\Z\8IW(d8:X:JJRV82Z/:IcLb:B/-[KDDgH6bQ
ZG0?H,QW^=;T##?HJCZEe[5D/bWSSd4\,/48B8<E1,0Ig]FLaN),OdU7#Q6U(@JF
</@_E@4A()9b.OVP-5bM,I,TUGF]SH6@/Y3<KAJ7U(W1LaBM9SY3R1]&+SU</\fX
V5RTD,fZ.fQ]=52XI87,?<4?GQOZW>G+[&5BV4UN4^^0\GW4_K&dDb]TRE5I)?aR
^_O7f4^JfBVH9<@2>gd&d7b,Ab-5PQ[\-GKR(0V>H.5</a/-O,LR\>LSJ;R0?8=6
]\FM6GSNL0Y:=8^,<)5&<1:=g]]fdfbS@eZ>D59e0136=4[F?>e^SQU_M4G1SU&K
=4?ZIaJcLaJX<#1CST?/?7+AbV2Ga9=,b_@-2I?5@:I)T-9d[<BRF-KQYe1<2cGX
Q\cf8D0&@D1V6F0.90;b,bS1NCbb==fc&B<DFFF5aNGE-cCY?M.1(b8ZF1>RFGF\
8U\cX\aZ5:)SIgZC_aTADRM5Y&&2V_:;NaW#=YZ>@/YQWTTFN1d(572GPCM35(6]
I/,0HA@A1Y:)]Q4+^YO=6@.Mg.V9NI;D3E^b4M(V\8Q#Q]dYVS+]DI/E58:A6]2e
J)V>243Q6]G?_;44V3f1U90dXVcaS)2KV&YG1[24cS<51Zg0,<>U+I:FJ:\]EfYP
UcCS3UX?.SJ4:JB?HQTd-G9.f+^QW7:CV<g5.YE0M>QKP(0[7/C/:],?6+D34&.X
We5-]ZBgBTLX(f;/\6H)?-JLMc:&Y?)8KNVJag6^gA=b7#LfV,FWW<LOGX4/OI?-
P^I^?VX_8ACg-35c+[A<;6SgOA;cSZ3ZACISVfgKZ\Jd+,61f=,JK+MC:OX?FVb+
Q[/dM:UB)]8@K/c\bVQ3HcM,)>:406+LWcK546_V[NO+10P]e0a:VS@1:[S&-PAY
3&IGM52YU0[Ta1HfIKF\Ld_UXLYb-PM8#<+CeE3GTAHW+gb<[dX[fI=]-cd6M53\
_+&4FJ5#/A[MVNXFG=a<,I91?1]U=1QZ;KAC\47Lf+;A=R6.R,f.UOfLJc+F8(&D
/Xc^@/aNMK&AM)0(PK\>/B#=31OS;GRaa/JY<DGH/[MC;C\,73&7LZ3dZCO<7:N?
b?6__BOX_<(H3H1\G=6c3S\LfF](^fb#aP_9TATF&9RA9Ya.++EF8#WPW/B,3S;=
CceV1N&d]1&9ENIJ8HH2_J;=J=&>/+5_GcG15ID?(35;<AA24K/eNA^K<>[M9b62
G[3ASIU7LS@=)W,+3S2gJCGHT5d^6Hba);MKc?493Q.87LDMNBMBb4.+JV1NQ^d:
,.(NNcWA;:B)+,V]cH^_eJR\Q,\A[,a[9fW8bO?M??PIT2@X-2(2I88CAD@,#K#0
CN#_X:a1S^\UM6cD0_UCX@2,U]L\/JL6(7<2&-714[.G?Fd#S+IZg0d11K(+^f;]
L_L^XPAEf1]]R<=eg-1T4A0KT7)+XH<C0XO:GHKQNeFOV7Q=64QG2WYWZSVb=bYa
DIGNN\Zcg3U_<.CCMNM#Fd./<^N/<Cb1.7R_HP3_-U,0Z)]4cJ:X]F)L=@cZ\>OC
eQ#g9ReEdFgCFH6Ja@b:d&N71<_;&3OZP@6=69:3d+XW39&Abc)#]SU_;,LGD2ID
g9?^C/20=_689]ZQ0BZ_EdK>7A#U4U4@-?Y5-([O-OP\4<gaZG.N-67>=a8Y-1&2
d;2P(.3E?bT3X);1F-QAQY;8?5/?[Yd-d/MRV]eK2>AFP+9D;O3b]b?ab4G^60L9
9\ZT-e,19VFeCX32?HfU1O\,-Z]>U.MJ_Kb[938&VS<J_-+4-a75RcI_@##><-DD
EKF:V.04+HNd\b>HBOR(8)JKWG^HQ;/4dB.c5b5KROCd6H3OGWPf+N)=6(3E+eX=
[TR&TKa#=B[bRH3Z,=0<-UO,KO,M_AfI5OTZfBX?LE,F+U4T)A=WcQKZ;.:SeJE)
Z\>HYa-g_AgaY4>Zaf3XM]e)=-Z9gV;7H6[6YIF3GD@L5L(fJ&FHWTCFZ/IBPcF3
WCDI6)d0EabR,,M7DU^RN8BcIG^JCT+NZP7;Kg\FFd)T6[0+:f]NNN[[7b+X02Qf
(W@#CTYBQ@]R134_)\P4=^C2TK\;WCUg02CTB66;2Gb5f<-=Q0U0W6K-.R8((79f
>UADI?--D=Bd+-gMC.eeJ1,gMRf?V=L#&fbdAR4&ENd)YI#V130N-5,@N7]=#(Z<
_fBDV^42N@fIGgZSeL>@I@Y@]Q5#:f)PV(b26/.EFX0AeY<_)9b8^#a]D^5\5N<L
@]cd0BX]#JUM0,./EE&OZ+P_NeGNa/I72cU?,AaZ\15Ff=H3<UVXR5S:<?^N_=Re
O2M\?QIF@]K9,dE,NZC/N,:WFaG76V\S18L@e9ggE)c2;8d-g/.gBFJT5>X/WYa4
S-+/+4E+?=<[#D58ZQ[eW/G5BHOSX^G)NIX.bRWF54]R3G9#ZT,+VSWgWSCMBP(,
L8SE-_888R/[)PN1ETUY/><26C:Y;U.JU7QCc\,9/1afX@<[6J2GC>Xf)A6+e)-H
>ND(QJfX&C@5E2S6&5GMV9C?d&3WQWd]7,,b6QXZB#HP_CeWPLT<SEZ1AB5L4R=E
U28KY;:J:=)Y,,d(LH3/_[6U[O#H#d^:,O(&MS>2R]1\#dXeY7bSX^0C0FRU8D.2
KAKN6__<XTY6>7;XOR>)F+1fM6I[S)FCE\@.DX60Z,2][9-6-,Bb#cR/YB5J)>BX
O?@G,fI:[bJE+PN:TV6?Y0.&UbR9G2YI6;5SA^cW&X;)eV&SIRK/@cJLcSEgE4Zc
9/1\EbGV(287+Vb^4U211MF<]P\=e4CURLST)ISb0/)63Y)S=M\RND&Ub]^1,2O6
<(B>O61eFJ+^B^01aZ:[X/BULI.7WK;C)HFfO+M87]c_?>dS6@F>;W/\B[T_C\X7
)(DC41B_8&-Tb/X_#PJK#:&^S^R6QgWAFP^UNFN?1Wg)=a(21MU.[Z0(.YaXQ8J9
_08L#9YUF/,0?)Z+27@90FN.KWe=&]_0:a8MU_@ZaX0E9gJ8Kd(eE(7+H\Xg9#Z4
9#6AA8MGGaIQSISFdAM5SVRe8L58<KG1_aSZ2AXC:J<a#OX6-&0FL7PZP<^NPUaW
C22?CSSQ;IY4<75<X#:+2K\d?Nd1Z^GOGdO&2PF6#<_OT/RXWBE4Y-PRHDa1EUdM
/3H_KJ642+H\IG>cU,M1SXD[X,I1T<?#(0C@Td(X\^bW;)QT_U7=be/SZHJDNLK^
@:5(_e#A;-R6)c8T,f89GcGA_7CR75(GPS:/T0=]X3#5a\d35DZ[5UH(9:g8/aKZ
fge,C>W27e)6&,L-^[I9.DI)9XLT.5(@HaM:D(+aY8E^\XA,7F?=EZZG@O1^(6Fb
SAQ1BLGE2//Hbg>-/4eH:02?SGVO.a-_\A#CI9)S(=]8g2/;+[IM9a7a6&X;-,9T
A+NEd_JMae74=Y9D/U8?:4@@@H#5DBM62?U8T)T=cC#g^6cc3:W>XMX:01FI]HT(
f;L-]H^1I-?,X5S9_a?9c>TRS2B0bcN9Q4ed;J_1A+W25,.\6OET#;O8S--(fEKG
DM\TTa)/a@RfOCXRZ@Z/OQ-N]&VTP1IMFg=81SIF8U4L;5K;/:HWcJV[?bVI/=OZ
e77A3C872ZeL4R7LY)B\,W()I;OdGRcZXEDKP4gVd6N/D;E2QKCNGC_=1>L/0@AO
;:(QA6#gYWXW#abEW0KQ+=gP;\\d6_B(6:5U4JY7R^EV\BfGZC>S4KY<CTJ(\f5>
V+a/a^TD1SXO?;+DI,,NXA]SBSXP^8L8#]bHZKAX7f-2ObP2b_-geFZ^)G/a-2WZ
P4(/)3#,^U<2D;^Ub6dRT+,+AdM=f\0C&(O/[9JfV;7;0<K;H:Eg#:@E(@>:B.aP
b<28#+S0I81eGP>JXMe<+LWCeB><1g>;:,(Pgd@6b^Q4_5KU^6C&0&2RV\?S=--0
CO>6@7/^@IC[MZ542Y\^8\W_2=#A.IFDJ?b&OLA;.]>DX/+L6fC3f:fSX]YH=Z&-
>T:]\\XFF1X75A-@:,1;9aOUQ;_0eQ1HUW:D@;_S][TH2?YQ:0CLKLO\NV-Y9[_L
1OLSKbNEF0;PP+TgUSFBTW88J:LRBGVbX>E=g&06,UcWKA,B495ZSe/0_TAC;8\^
].K>SM=SCQWQZRaIC3,<_(2V&6f];W]L<6cF1NP=W;HD[=6=?1^,QQfDFKEG^KCH
4d9OBR+gIagRA<_C9,)41.8_QW\<fDF&FHdI6_&4+>eW<fY=8))e.8]W_N6;1:H@
)Zc(<\bK6@2PNEV;\+TA,E6Zb.9]G5e7RNEH<IS+5=6/2gZQ51=52d01fU>NaZXa
XAPVdSaP+/5&FC8^2#P1^JGSO:QTHc3Xb@Y.J=Z.&F+15V:?Sc5=X#a-aL\DYJJL
_?-R@BN[[fGfK^dF[TBU)ASY#gUKJ83UXE6GW6@F;:_K9Z3bZ]f7-@IVR,,gR:9\
51>F6J35U5(dSIY=LN:H#>LMfC@eg7W:>8OI)1<VO>X,;bVaM>8\aacKBXWLB?9S
-0[SSOLCgZ\3CcM-bXN;8?1fD=ZSBCTP&<MLP1VK<F(^3=.GV?2)VHMI4YEN?3I-
<beZK_Hf_DGOaA3<T)95S;UJ)YC7ACD2#6_;BH7(T&eRS<2[C>I+X5^e,LO6D#.2
(2d2Xc?:&=(54IY&7U,c)YBGS#GZ(1M,\:164\e0&5JC#&39;-cdG&<YGY@&[L@4
:25O_)O>IPT8^V4+V?T@b2M]AbWeZ/B):gT<\P#+.1^1E^H#H-7>W^3;QQ^@(-7c
Q8VdG[HL4<dJ<8AG)LNg</JX&N^5;8)W<d)3a#=HQS&L/(I:<N/E3YR1AO9;CO2<
G\GFPcHH^;/70De)=V;eVW7bAXT:B=6-VB<@,#L?#WfNV])6/1U(HRf5QQ9S&9(;
.,ddXIAJD/W60ZY,2B297d)7XBXH<I40g5dLW19?3&NF//[6ZFe(T<A<6e^06,3H
2Z\QZ]R7O@\5Q]g^)SbFQ4MPDP7c1#@((@E@Z-aEbD\c=/R(d94=^WbCB#deO-JV
MeY+/\JO_KMHN:CQ7,XAF/HL?[HZg_K6;gF6S.QFF?78BM^85S./KRH<N-^cUF2I
+5P1g70.88[\:BZT6J7b_](_PA#SOFVIYcW@&F7-FUS2;T,2c;1B@83^&6,QFc4-
V+d5.ZLFE@(#1LSe0_HQWNG,aR?B[_>NFPbQ4302fG>-3MAc)4(OZO4(acUVPQ=L
HDLbG(Sd-RYH\#@H-KH;F-1O<G.I^JB7A+A)4T)c)]DRCgEP.DGAVXW\-eJ\U7\)
6+3YC\1cbX\Ue&:dPcTEXbcfKQ8dQD5?C403SAMPKM_cAdAM?@##H\&AQPPDW(YP
:W)3Y8/>Z\UKC1<WYY0eB(&Hg<\M/)CYC4e<_;:>F3HLfSX+5NbP/9&ICJA?3[f_
4J]-c->U&3L1:GIC,.V\SdgF,_D(28YX<aH#aMG>K2E]+ZTG8R4V#/,77RZNA@6V
a\aKgU-_KH.&CK=eVc:9CU5b7R/K3\0K8&WG^80@6]Z.dg:Q.\V<Y86]2:Db#e]1
3XT9F1&<3NfF,-@(?AbU2=baLO#1P2YD-=WWAg3?-;FF42a<#.M#ZSEQ#<#FHCWT
TG9[[YE+MGI6fR^>eP.U]bX20E9Ga&;Wa/MVO#E]X8bI>W<4+g;3>&d_UdK\]R)W
/M]V2[1^[1,[\,JTgMD_c0Je@5B6Z--4@aI@W:CPHgN6GBg1Y?T@CdJH+OS]9)bf
8/7>8bWEL20/@[:B8:8B,FcCVc=-C7F:(d&O;cV@VDH^Q7G2T@ec0?KON:95F.-#
[e6F-B:7XSg@5A(]7:Q&D=Cd6,DCL+Wa(^/ON>&0>GWSU1c_MU[<LNNTC;S?YA=f
GTUTU5:dIE3>9\=<&LT9P7a=P\6Jd?H;\[1DEKb42NN/6+&b0PIR\?<E3C?[WW;;
&g9CeF1)NCcGSdG>70.L]EUOZR>#f&W.\?&b,COd_:)8NHXL&b1:8[[>(+RbP[T.
]0HB6?4@5f<_M4A][),QGQJIbFPB1P+YSL<(,+0^0+V,&=7L0\]g?(1>T,ZH#D\Y
_7g)8Y@^aAbeU@S<+P@B([FbX[7OR3_S_.FBY)cD?3Q3Ca8/P83@J^WRQ&FV2GK=
8N)dg.EFT8KU8^4#fgHY[O+)IF/.)BW1(><KeSSCS23,^A^T61#.(FSde<DaDcKc
?MVX[D\KP?QVIcBfH+O_<H<O[ZKZRA&5?,,KKGFGOZ?8HRA[5LM+R93NCc;ZHAGB
2Q\>IQM8Y616XS^7>AO]E/N.&8;_GPW5BFUc3WTf/F8d#[Jd:FU;,X[\?@K1bZed
CPT+KX3[SeE_cJ.2E@@KD/8//CFG=QV\,O3fKAJ:DB/,Eb4-BU37c(4cX.T](#0\
^P^>Wggb@FN,PW^,SC#0WJC?C4d7OeETA?Z7,6U-M=5J8J?JRE#LQ5J[8X1&_JKf
R[,/8Ae2G+4cIgOXKa@-T92d^4.2R[QBFcDf.QZ083@d6A/c<e](AV[EG;A4@eI?
b<dBBeAPH=WDRNR,a+.A3#[D2B@?OF-FfVYb&L^EO89AOe4,4].f966PgWa-S4\#
3bf+C[Id=/D3QCFN32@^0VC([LffXZa,2f2AN^/U0,ZUENV#A9U8)D<?^+8RYDDf
eDeDX4J=_f<\Y^?K-6B[1<,PD12f@?()9fXBQ[LKPQ@C/531a,US7EEG4WI+IPcb
ga>J.Q\2cR3\(YS1J?RW-P=2E^L09]BE>eEg;HJE=7>6Ff^Xd-6_GG3.M>6LTRXW
[+#(<)eK\NH0]T/S\MI-+Hd&ZNWC7FCMceL[K<^QGa1&DP_##S3V9dMQANA^&=;T
2ZWW?=;fZ<#(75>M^b_S.bD72MSV>??1c.;8g/LTD^8AeFCB/H>C]N4+1QSP>b-I
\3WWN;+.Aa86ZMa=>?Y_RRH\7V,Z6a@Ef091P?f;FKZ(b.]+Q:V2;CX:(D(WDW0B
LYRe)ZVe[=A^gb+SM4/BT&HG@VXg[ZMDVa41DZ6]T_11^;4gA1Z9O>QKKRRb-YV0
Z>WGCgT_^W7KRLXP+D<Aaf0^.;/d5>>S91(@OLO&3_b2S,F4L#YJ?6WF.7L]&3D-
>E<<e5>PJ97K6C=DAf(,c),b^VE1QLBOZYYBM#^W&=[1#1gFJJ8fJF1NUc-U+V4X
/\5ARN?Nd?F2a([H&3/W.C^eSH72AMdJHb7;bX<A+^ZeZ1J.CWOS^;eD85LCdAS?
S3GX1>A#92J;&Y&cRA2\IQ93V\S:^N)1R^8&I=),Z)1X?<Me:bc>Ge_0[12<YfAP
CCCfGf?</PW>SIWb&<0bX=FXf/R(e<,(<8PX=Eb<2[+]V0,00K8FEgf:[(\S##&A
dH3:>)M+5/N-?UbQ^@]5K(LO^ef0Q,GSK4d/SP)U>3.g&9^.Fed@.8-FKFQ\eU[d
fcO<FK9d4CRP^EGA4cAIcbW,,\@W@\1VR;5YJU^a?KRTHU/R#:Z/X@T)]DTRXL<W
03/g9U&Za/(HV+W)HFE-H?CIVLCBeFBTK;TTVQ:E+Q9[]@_FEU2Md(VaK8BA9\-R
?[Ifb/ZHIfeQ[@)7-a?UFIG_DMc^.=N;HE>d_C(DFa@\2(8/@4@KJ1D9)&X#4Y>f
BaT4S,QScJBJ0;&C<+).fAZdFgI?3A?beR:^OZ0[DT,(V=^<b@+X_2c^/Q0,Nbd>
3YA-g:<eb12&a+HWBZKV2G2ROP)aI1RH&/A9L[]2Eb,cbR+&G&NNZGRB>#1#]<a=
LBfCT&HM5SHIfF9H&B[b;YeL+2P^B=>^X+A2(&;g<?=3CZ:cfZX#8/8(ZP7?cO@S
L6UK@J(D@Sg+I7,:4-OJbC\N_ML=b8<&P73cX4RQWe_?YUNW[XA.FcF;6WI<X6N]
0.H55&:_a0G(&VD\,#\e#WT=)HF-/#8(TF]P),OW</WLMITH^8K.^STH##dcDH+a
Z?I@b73eee7<8A9GB3+F:IbT)7E(>:@=R:<G\Yf5<[f1O_Z#@6^Rf/LE]8\&c?.E
=f_LVO9fV1@c\7.MX>eNSL/Xc6K51[NaV0aJOX.E?U+Y+AF;<Q[B9<+-Fe.F_YXP
U_8ZK[?\+GA8Y,040MT6ZQb+0-P>=W^cZN>MK9\R0V\(Md9LRc,/@D2b)A,B_e?^
VFNV5SXVcM&3I<GP[A\0HJ@_@S0Def_TB_7b,aC4LF5@.?&-G?>,NK>SQ;bM8g\&
NfDN_PK;\4&Ae)_dT(cEVJ\LNVHUEGZ1PgBd;_?LeYCK.5]I46^)]M2.I>WRNG\=
+JF+HR>(bQ8548IY;/TBA[f0A6#BdJG-CP(M7cb)XGc=P(2C=dF&G[32/a3Ida=^
,d-7.g9(2._3@K(F,R?\U6bYMWZ34_?R(a7F3F>[BWE-;([Bb/H]<+BL0dYYGLN0
66d+Z+9CR=7F?ASa05@R:+O^F+.3Lg.^X@CB&KN_E.G4)0^W@]S8.->7KKSQGKJK
&IXD7WD3Ee=2J=MNB2Y3LM\UYC.a71^]2QG+V/QPYK_ADEBU\P:FZM@IHgd2#O.0
0;YC(ZHT2_=f^.ce=-]N0[H/E8T:)P&e^-LNb_#^AJCcPHOU7E>UNS\cf=9FT:g3
Pg0U?9P7BBQL)(7-Gd4?GV+3S7c=HF7@0\0]?1TBOC=6HC6VcSNBb,#<dM2ALf]6
fH5=:DVd[,V:-6-)_ENWW>>H9\VD,Y[EaK#\cJ-cd)Ggd.;P.O(VRL=6&d1VJ9]T
P307GdeT.LdHA/G.H&NM+g([W)F=-g@9EZK[eJA5L9]VEcaQ;/7:7=3>=7WR>-<_
#0BP7[(5#(U=d(HY30)0N8X(cQ2fY5ABM>OJ0FdG.=4GMLG91<]EIVDFY4:9@[B^
,ZDb3M;^TH-ed@U[=6eKIY2.3K0W8ACKd?\bQMJ5B97T)G#RJWPNaYC:(TEa+I:1
DK41D3QDDQdC)gTXWS&HIfNbB)eb4#RBH/EbPg3NPUOPR^A?>H=(gL(O-gA\WU90
B1<I<aR(/J(V</_a4S#622<Ibfb48F^6]2;C7agG_V_.cJGcMa&+OKB/_GW1^E[2
c15/\..A/#X+W[R78;Q;5SK5Q53G3R:I2&7BOV75bO]?N53gOV;WY2eZAUXCKY4>
:ARJ&_?IJO&+cDG270&&_C^L6(bNd8@G39-L6H)cUZ6[c4V70]6N@ISN79UENI7+
EU]?S0U8PIZV9H5^T)DN#F]T&\DgXCTdDbET^2R#S5;Vcg>2PA<[SR,GT:E(#3;c
[JA:g8GBUM<T[BGGI4-[M,CFD\eYJJ5QU(WB9T996AN\QGBL[V12JNK0aSOILPBM
(HB1#NKBT8gUa(]Y=OUJA\JZA<(b0S0U#=.A6WaC__:QQ8TOA;9;aNJ=f/DWa(S#
6165,UPg7Y&8G=/MAD8\:KN:HZVH6VCZ>?8TBg]Z96H4QM:;:O)C&d1:>A0Ue>)-
XKNOf#BKDT4bY@dJA0X/E.P\R9(6e,IK]a7GB_BYZbL]3\HAfD)a0V;R7_8\b1(/
P]03P.5&>Ec@g5IYQNO0#OAAA4A:.a5F)VRd033@Fc#LN]>Z4:I2b(68]/.C39F2
,VCd=RR(3ZRX0=Wb5/URA#gRV8\>.H9I>H7#>9\6]+A<AfK)P)DG),V[C)e=Dd@B
<W&.eE(D,^[Og/]@R.gUJSY_+6>;(3;5fU&D&Y+QG@_):D67cfG8_)(<eDZD8]R-
E^4_YWgD]@VfdOK@UEBUEAe(.NOFFU7LJ_<R0>W9[;fT7I:[&4[cX)&[K>8<#PJX
8P#[=L?>K/T[<X9BS9ZMY\ERB[d.BG7>(<FWfcA?)Ad(/^7DI+#d2U\.]^;RgUO:
)B5-#?f2QM=;a;0RKZa+[_DWPF?<._97d)2EZS:1K:4;GG^FK-.OLf:f_<I,)?bT
\\5E@IdHI_/c9ZUXc\&Qb;?<XFY1dd<N>4L6bS-Z@XLUee^QPW_L[g0Z2eH,N_#Q
.dOdN5CC&^P>SOK0:>83UVX]?SJ>X?>807Ig,-6_OZ4?fQ7G<EAMR[<^BJ?2SJ)E
UT?fT1K(=&3d26R@a><ES;FITL-e-MNSgRJ.<7.@(@P2ENF\U_@;cabX]>#6P\#O
_>9Y1\d..R4BBJgG4NK57P]FM_FDE>91d/VcEZ)c37ISL)3&XZ;(TN(X7c\G]>cJ
W=YREP0G5cC>H\CUE+M[?_;W;UV:+P6=3<V6;NV;2<AT399<]ICP2,gUDeMM.A=d
@=^0@]a[=N[>\HJT^_=HBZ#>NXa_<f<G?@7\=^O0;]@)\^0^FRU1?:+,M3ZY^g\@
PR6NUX6M2(,2;6AA<0M,/UM\:&U_bZ\d8+J^/dO+:(=Q[+,0;K4MMYQD)88SZ55Z
SUgUKI&X<P7BW>@01H0+:Ta?)<RaHdO/7_PW3ZQK?.T1^MX1Q3X70.Ue:51R5PBf
4F<QcI^f4Z1bAdFX=1cQEX-:S-R622UTNNeA&A;_6#UM,If/^2[([6_-T1VJQ7VL
X2@J^8V#QP/Id-XA0<QO]R:+H@^3,YXEc1+OOL5Z<CPSE82>.^>^<4&H<a8:caEe
RU9)Ce9eGKg\TFGgYE9V_1?dUG95^Xd3A57ENE=N3Od\(N[R_/?5J0)_7a??9+T-
.UW?O3WC053T12;=EQ>=6F3);03_Z_cFc9PgU<,<R79bD6]2[<e/PRf3+JA[3F,#
N.2(C(a&1.dR@QF)X6,aN_UO^ANSOcP4_6ZINe]:A7KeRJbL2OS]3d?(I?UP//e\
U&^S^9W))JMD1IG2VL@DZCc(R\U45f+O@O,6_IHJJEBN:e)5=^1DQD55-,>#&\4f
[8C>>ZR6CMH-I/]#M;^O6Mb6X)Lf1>b/0GK&++T?.U-HQAMS,GB@W<;=YOO>16KM
)CAe..@K1B#><V6.Q5b<+(X?31<Q64#ZCC7)F631+-K&g:HMeXXT,J1BF4P]J9cg
dT]+L=[.</+\(I<9HfIG&<\3_VSB15VF^N2@YNXS098Pf/AGQ+@D2W_JY.aYQ[(1
;-+KN@,.\9eO-e>Z^;RECd9fPbC0)ERY7]Y;6QV.6-eU+V=0@EN06[BBHG<f>aM.
RKK[)TcBZ]J01gVS?EPB[NF,>UbgB^Y.UQ6^\0V[EI3,FMXFc)Be,)7U+b1:6;^7
#]]@0d,;-THKJ9(T)O[@0J=\LRUFO8gF+#0ab08-)\6A]\gB5Gc5\5XZfYFSVZ\b
,D4-3CS]Q\?c3M7_TIU1b0J4eV)_]ZVSV,WQ;GTULIG-M^Q::Q?X/e-:-e<(#2b;
E<]5V28)d^FEXY<O9ZXUQbM7I0@Fcg7e+_4[gb6=XMFOG1W?<&G9JVY7HV?^ZFDa
^C5Gg#7LB+TfFL7_-C3M?[[Uc+S]a59C3XH1G,[;=FRW[OCTNIPCG@daAfI4L:cW
-IZ/cJK(_I=#>_^CbS(OL&5EA+VW(#62(L?X00S?1a^93+X6T6377-fGWZ.98GEJ
_[(S>M-aY42Z(+02Ad#_>g;g?50N9U8>C]IT4JDJ4ag=A;4A>,OQd(+cCaCIHa]-
BeT6WDXb+>97W-)/,CAUI,6RHD?5cZ=:A>J9fgb(6R]Rd4^:I</<=PG9Gg>VI^-O
^.LA0eM\YKfYW#TUT^e4;N>aT7WK-fK3ZB(9][\E<4\fKP1HSKJ)1;RCXeKMXIIT
4b-Q_UZ7>W2C8^^ST,MPTe7T71LHdG]3D[0H(_bG(BNHaH4]WbH[^Y^L=F)IPRJ5
YU5OcVL51SMP?5>RR;,^_8V0NH4fF-@?GMA951T6;b7b;G6T-V_9T)a)ScX5be#P
4d,<gR?AK[7ON)+03B:..9Y8L#NS7Y(ZJF5ZZ(3/G3Re5R1#)(EgdFbZX:[[ScB0
#::79&;>O1N83\c^]BGX=fdg;;S]Ib/X-^Ybe#WI-XBVKM0D?FDa.31,.M<\WQL1
EUE7T1(0=7d^</7P?cIgCLg+G7FOKAO2cXQ.A=b]G^C/HDWP.\a4.C&V_/X[:g6G
GcU49R3.(dH@W\]a;3Y:CZ4?G5SZ4g(3WGC+1D/e]S[->NAR)7+3[?F4042R5]0V
aX&\M+(V=R;.D.b1@K@ScC])Qg;UHf<C@P4bb?f,5ZYX#AA,BGdF1I2&+(d::S[_
MGTc0,[I9dc8=^g&2<(C=31?8gTg&#e\KeaQ]&[g-af@LV<KM_@+7a]#0L7WIRT0
.1D\\_6>fSdHV+9>:gBJ),/33_RWP[U+/=OYBgHIgO^X1X5XY.;4D;=VV5e]PK1b
@6d)REegAd8O@&=[gWDWG^KdfP:0-N@X---?]A;9#<W-B;D<=)Tc6B&aM[PVH&-,
Z:ACW?XNU7W/eQ94V@Gc.BJH<4.VND4ETOA+Q<6]VX].4LFb.Z2gN0_X<E1ZBVdf
LMA]W#Z:,>e0dU\/.&A7X_DedS7N3\aNCVG[5VZGaaCbSOSZR9JHTd=,\e1J;_A+
[J<bWM03_c.7PPU.W^V/3J+W,g<L6J5=#(-Q:SS@Q\5.SVOM&W[Z,=,U8<P0/VJF
@ZE7I;Y19Q.fa?fM55b7@]fV44^^(4d8?D]HB9I&I,bYGI#EB[P9SKPXDCE.FXHg
ABZIF4L;HPe+ZK@:BS#?MfPb:W([Na(DQ)\gIeRMDKb+Q@UXY;QOWOTI-PEC^[d=
,).cO/gX6_MX<5d([J;GVPW1MF+5?/@4>[;g_[[HN1g?26&:.+3#ZOe;;4N:;QdE
;T1Rf;(bL66_FPTP)WdZff_XFT&;a\D2]V\]U_f6(:_T0bfH-=dH-K<[:-OL8.Q]
V;A<)+N&ZE(0>(]_<c5>/]3X7_W7#-66&]@M-b4MZDCdcYaB3ONUc@BdO0>GYSG]
7VRMFV_9V21STPBZcBD#\I\KK?c/fV6Q.0.7SZIYL1f6\P:N#(YSJK_PN?&#0J/D
=gNT,ef@1CYY?I8#=A32=Z+E<]=10GSC4)A^CaTcG]S-CP?4;+@BfDT3(A<QQPU<
3#fO.M7G93^FJ2C[5df<b:QP4bgT>df)B^;8:_1H-gK#)STOeO:8Q9DgE]<bK#B1
6YCXK(0#/&RO)PU,N=f?8B^Y35MK;-ReVS^Oee#fA,:8FPKJ3V0fPNA#U;9aKf;g
ZK)&I.06\NVd.7Q0;>)9ag+L5;F,?.SH_15)f#-PT10_TaIBRY/GH-Rb.Cf&gM;b
<T3Xb@H5[2XKY41PL7]5@MP2<56-2D1C1#\R+[#(441/R_J4/gB7_F(4\XH;#096
;AL2L6F6CUJYYd@/5/T.+-A;<e@X/[bJ&9.PXOC=-UFbM\Tff&6X?(#:CT[^)0WO
&#8A-\dMaK/7J[H5I#(4G\37(U6-C0\fPB><GbE=Td8Z#W[b(&0K]7)7XO8J5G9E
XgIBYL2aEQAHWF20:,f(1dT&I=1X9D_Z#7U=^RR7YTOGd?KVI6-4@?^,dPZK_g/<
ECZQDD#X5L0KST/EW,e[A3ZA#G<FR6OXYU75M7LQP5C0/V-g.6UXc)P?VSE46fR@
R)2^V:;If=:_.\>ZD4e4;0>MC.##g?b5U.40Ibd9Pbf[UINH2O].4EbLD/-8BYYA
]DXPTH^GNaaS:5fe>E2^c<,R:7IPPX93.<bW[U_YJ(DTET,T1HSSe,8@g;@RL0RC
FfWWXLV0,H@6YG)PHF@,TTVWR_0DML4HACH375=^)cV/>\B\=V7TbBN/8-ALM[B)
\,QHL_E.+N<W)8f,S2H_B4-(g#eKG1gf^(.&G.W4S4?EK+JgC1XY3fP:R4^bdD4^
)6\VBA3.0U^ffO60^dNA(22OU,[e+d;LEHLW4;7:93]<@95dDR,5(P.A?9gRcI-E
1_ZAB/3KOe+.3)?8/9S=e,34+)Q)>c9.(.21+@V0MVQ/,bM54cK7:W6+]@IB@_?.
e_D9&^1bKeR;c);.+?0/(3463/JE^].\Z#PSg&b5a^0d,F/GaNIggE5T;aYFd(FP
eT7X+EcIP],P^G_a?A?I:.-#W,,5E1Qf4UDH4=Q0XFE+Ng846NANMQY6Y55N;Bfe
S96g18g-\/IbaGIRW>?bAP1G&0_EZRHF?8+b,W+PCXMd5KO2bP[/L=0T730LfE?H
@U\>1\WPAb6,;/BNK:b6.D<RLPHG-&F<XTC1-)7.7NE74KABT6bA:8^(fY\KcKe]
LN.O5[\-?X+8TY&SA52[@/=0Pbg]AFg7AbHKeK#]+=.XFZ.;8(gJO_CYdR#a:PSA
X7_)d\?bXO0=&TK6&dW,+D[D2ZO]J;L6(7ZQ39S+PH-5,C=XOd/]NXGd67S2cB&I
EK:cA/<fZg?=;Z96D.S1-D\cOBaPA6?df/06/f-Zd=g&B)J-OW>I?3U:&dFKLZ;E
AQCYWTZPH(GEQ],4AVbB<62TMW6aLSF[L0&S6QM3MJ#8^-JX(O7+7W.?_\7B&440
RY;E92dg9Y#6X(cZ.)#F\g:CK[YcccWHT?7,N.]FQHb[X&Agc3/N>G@N_B/e^=EM
H+1.)^W2IIDU[^R-7-=W#:U5-+AN+P-+KQGMU?\EMRe6;G[@<)44SWg81bd>@U/a
2S#\5/VOOI]ZCCfJ;P1G;L\;3O>C8Z;^X7WQ>[Y8.B9eL&976;#XX972g0&IG5>1
(TXXPf[>^;U;Z#?TJ@(X^)2ACc?ES>Y6R?FaF_IIf4#VSV;T&9AA?;Y-[01,g[1I
SL@>eI5QHVEW.<a=:SJ+T[9O81A<aKXb5_C90bbdX>\d.5:IfX#_SQFJOUHOee]H
Qb(NW:=a8GO-7:R.H.A9dc330_ZT9(\]_95BCdVHE3QcWI+3521,W(\D0K47>OHG
A4_#g[P4AfJTSM#^V,M=VPQ5RaKfS,YV387CJ\Le^\_^XabKTD]ZC3;Q><ebRZ>T
7].P#S8\O,8T3_TWF6?&KT;=PJ<0:13(b#_VXe\A187[(Y>@0FM?,7Q^_@=,._;=
HfS#I;DH#dI=IKP68(K.c(b2f/4NJLMf5W>585be4PY,eVTg/?HFCd\dFd,6;-:R
c^VNdE&5.=.-UA;e<2@8=OGQ2);CKOX2Iba71Udf2:ZH&OT^9P\LcB1;1(FH=JY=
T]gfe-[Y#.CH_<b_QF9@IZb@:GW)]VLY8c<APW/Ze3Q7;5M4G.L03a=);VeXR_<E
95>g?UA,3WJdcG\d0U=b<9O-R0BNFQK=<T#H+&RVOA:UH&XX4IOeN8DIb,+VZ1F-
#VZEdNH4RZHOZ5NV<(g;d\d-e@aHPGYB5#?RT-7Tb8Kf+JER]^991B7UVYb:30e/
(HKOVa^bA-&20[VOX+_FcM6-F+(-e;[ab7:-E0-=Ha3YFTUK0LUEg#Q,P[Z\WFUP
A.57O&)aAZ5g9FBdT3P<)e]cH8L._W&45.=5SV7W6TKAU-[dE_Qb:8VR8(#O]=PR
QLXe<[N2]\@OU4b7cSR6?3fR<]K@Y:.8@+(^B@Z30F02f4/WPQNGN\M_Vf.LS)ZZ
\]SRNgAD[BL]6c&FN4\HIQ0^dM;dC)S\Z6a/>?gGINMa8&,C,>HM5ac8V/BMP\DM
4a/@9,<dG>HF4R1.Y;GTHOY-F=^O[OP;#;HF\dLXB(?>I/QX[OGAfBPMWC:gO=JH
ca(_5AWCIDR6OX[aMPK@,,b<S-_I7WV6Hb6>Z0(]-+G:G\SdH#>SF@O/EBd@S@0Z
F,eV7(;LGM4bYW;>NgTR[K(QPQSXdZ^_K1T=6A)2>f>DbL4&S^WKKH)4f7c?)AZ9
WUggR;/J+(G\1O?,NN<-MM=OKZD3,6WOS,Ga9C+-d,@cO7#>M71N65\N=4@G\(\@
FeHQ:fQ_BEb1NUV3a-cH\Be^0Kb3<,<QZS\5C(B00YAAg#E84eD=;bee8EJ=[b<7
cP9>ZJFLJFY>_Z52ZF+YJC.#51YMZPQI2b0^]f#+gJ)D1/I+S;@.^3+\IJ_]H6J<
;0N9EALV.M^+T)]gKUV+UU:S&B?gX;/FX+FNSZ?B>f@E-3KJY&g-76@BVEOGfAXB
O0a_/eNTe[^/b&ZMY6>,:c,J0dbb1]Rd1BO&S9eQB-_L[^L/bMdM#,,&GUL^#T=]
==FTb<fb[Xg[@dg0OF7]0;d>LO5<B#.38J42Z#6_BN)aP>R^NUF.WRDBW>.?c6Xc
6416RL\bXNcGYHRV;cWY\KIg;>V;,^,U)I-.;]:@]Ie(.VM;9/<ZANEe51Qb#-aP
]PW5?^7P3V\7EBXf5/0Z8G#I:PO>[>HcV^^,=+W#;d8NC0AR@g]4P#JJJQ@M#.;+
0XVKG&.XQg0<]P[&F10./;CB;<&+/cME?0#/Y=ZPWIWB^(Z;c0]LP2(ZU#&Qa3UQ
?>f<@,c/\XZ\T_-PeM9C?F-APY@aN^gI6L7BEW);Sf_g_+N>JLN:1F-S0bE^-Y:)
5;<?ZTCY?X@UJC=0bZDfa3V4//8WYe97FXba=69WdX_>aa6JB,Q:V9:+C1KVBegQ
X<(9Bc#PT9I@<<Ta-P^S8ITMV=JSUCaU#f__MM@&BU;;,7aeQ6&&2IVPaI.@G5GE
04FB)HJYHU11gcaPN40LRa[P1OF6T;c9G+VX/.MRFLY&QH6^PPA4,.^LLY]I</[]
[,DdYR&=2gG&-J0S4g^4-G/>+ZU&ac2FMA5SB=<I1,bfV^K1@PR_8B>ZH0WbQcd8
A3J>a1VC9UdESA)O3-)TEXCBfb7/FFdbg>J38T4dQ22ZL;68TE([O/FgU2B8=(;:
^7@8-4If=AV6SD(5(WD+=_Z0&TVFIAb15DaTW<<VNWL[?9T/<];(U/d35P#]<(JS
:E8//2Gf<3Y^=^dF6ADeLYWg?HSJ=;SU,beN+N/#34K3-10\KDJUW,-0>XO>]bL(
-]<?L<OfS>)F;GSI476_E_GZCXdE[Rf5NRFZ>>H0eYd;D4QGYaH>0gY0L89:^K1T
K=KE.O8B75Fba9>[+5@E&>4,bbN1YNELLM:R1R+\K5N>Wg_+;)ICfA8&+TT3,IJT
LgIc4[V:=[/GT+BE>@[T/_Z.JP4MO3G9O(YL5;ML:4@QaC]Ne?HP\>U31e3[M.R[
DH1P^-@&Ad2^_0-1LY+Y:QQee9eR786)D73Y<5-;_S(@2\=,SAS\[.&/_e&4MSTf
OO9<f_NM?5W/FQKEU&Y?cg6JQQfI<C,&8MB<&=9X#g&0F)(Z-7&9dHIc0652>agd
LR:W@;Oe#fFIMc_ZW9[UXD7#.G4H,(B#^2&8L3=VAX5N/MZPH-,G=KJG<2QR/_)d
c+\ge1d&MgDMN:0<=C#NOHNF]a7L;O1c__?<W26U#R[UD82SM>?]U.:[=DULU=9G
&f(?LCg)U8OP>[W25b;Q[R.4d;XELbC.29GBMQ6bfP41/dKNZ8IT.F2e^:YY0cVb
_D1VA8MX#dVVJB5f=<8a>?F8@&0&@fbO05?C(D=d^(#\AS(+5FT-?^CdI73HJ#C.
/I&</7+H-8L<^b-N2)U+OE^5,EPb8@Be(PH.=1.2G9gST_&:ecHR(0KY0NVQfA)=
SQL=@+-9D2f)VY2=WY@,<Z/&N]:^HI/NgU4Y785(@WU[VM09GKYdba7fIB7PfF?P
JcJeBM-8,.YB-G4[#TL]5#?f</-4EMUWc=CFQJGF12Z;1;B79JFL]C\P;?b8(2,X
_22Y=1]-V9^F+Q&g[5;MB/_,T)/AUD,Z=MDP[=[e\9;UbA1MMc;&\gT2[^I_bDML
\Lf8Mb[3;L/Qg])FdFaSE7XHH#Ae7:KO,g247b8<f:NH\O2(A+<_d^V<U)TfKX0R
8N(P9VBa:)g]c);&\[PN=b:FJ5#@((<G\X]828bcU^adFJE9J>^=NJNL)&-IRQUV
XH.SPUET>TXRC?X^_14RA<.<B/F.+?OC#cZ[Vef&;A2gOOe16Y<M-aCB:RRAA^46
X@7K_E+]-g+=./]RP,5B\[\Y@WUfe7]G)\U;b6U/0T]f-&9.8<@C^7,fKfUFH61R
g_-7,C8[YUFeIdSWE+\7e2/O3,N>I^A/.AG#aOWV5&?S6A,&LOB(Kc84GXW_0B)T
;;N#,L?^Z6d?CE,W=QA1BZeBJ(5JZ41O[-ZaEc)@QX4]51E0/d2a&SSCA,JL4fF=
,7[>PCH?IML0<X3>0J5^/b[?Y;Z\,U?TUXB\,b3&MBW&TYNGI=5+#8>[N@3(aV^X
Xd82OF9#>X5\8,\a?,]#CN-ODVgUPP)M<Y^7TeZedf(PTa0He:bK&&4?IeV+QSE7
73YUMO6;IX=PPG0b_0]L4+64,d+bL22(;)+JHSFAK;&e8KB\ALIJ3XR3(c,O,Dd2
-]GGgd;GKVMM2eEb#<P?X#?)JH1.F1\VM[6Se<Zc_L/g,)NdL^4RRb7[1:@4,?OW
EZC@=MY-KJ^3,Q3Y+_A4I[SIaC:/eZ=6eeUGaS.8EXac]:D@<<+2P9:.2_e](c_#
.S&NbFY&If5BSW0Z[(?TS.C0=R:RYR9K,3=gNGRAfV\#V+]5)I5Z5^aH<GZ0aBZ/
[[Ed]U>+NTB(A^^(f??=RfQIZ9Dfg^LT&4fR#7NR0J5),/8A8G-+-0\Z)Z2G;Y\P
N)HZXTF&<=C-b?TQ9g?:=3EDGS.1BWCc:ACZ0C49;eOXMC[VBdD1,,N<]TO:38d6
SAQg=:W3IKN?C,\H]V@K@Ff9/dA_YL8Z2F9g2.;gB+@(U#\[=Y?6+TTY/eZ8V@O=
__O:W3L)5>N\=IP7OD<UE]f?]4#c-BO>=7KTY#>&@QF963cOdY[DFF&YINQ,B8FR
AIVeOabY_[D?QRFbBKWcY_H>6.]R-.I58TfRHVb[X4\PA;.44[A:OgfSB4d5H3&W
=]6^,-<6JO[:Z7L2D4PI5WMINNE9^=:_PW+-a9ea6V5RH8V_L:8N-7GJ<U(P3<.)
K)A5BA=^TSWM.UdXFM.4)J60?OOa^-[_<NAQeYH4IdX6I_Y&YM]a2X6P[14gI,9A
aEW?VR7fe=]aFa5B1NJ-?W->.,NJedX+cIf_;g/:<PR5LTW<@Rg(d4/)f6\#DeM.
3?WZICJU0EcA^I/JgZ@>.MgE9a;#V0X-=I&?(:2M#EV=O#A>OHJ@ae^de.Q^1EUb
[KQ.RgFgQZ;<H9/eH(EPH>2=1]FX^I8+^EQc/OP1UZQ2H.QZYD8ZCZXZYdeKc,?T
afe5CgMY8JE&\5A34SBA0AQ;KZ82P-8=)L]a@,d:<0/^EHY3;X,^K-AMVC?dA7TJ
UQf&JfPU5&[-I+?gB-8/^A9?dWO3C9G79-6cYa[L[Cf[D1WB)A@EP+[cSI:H.8^&
,+FNNXEX>&QH4_BKNeZ/X;4dQ/^Z,]e,2H_I#[NVJ;;Y_CP+JYbLZ^6Hc,/S]@b)
CdXX7=,2:-?:C1(TZe?=AK7_B\3<Z4_A@(X&dSL2+.0dM&,I+,JQ@YKFg/1TbM+P
N<<F55_,95H1/B[,^ZeeEB+<,X+0Qd@7gCR?daEX(OIEI#d:CYd393LfTL_5Y8=J
27Z6];S^SK@9;W.>b(K0Q1E(cB(4R&)<ZE,00XC297_,U#bU?<_fO8b(8@9OgVTd
#fG1491f]I[KXb./OR:P=V^-TOIZB.[Sg8(.39-f7Obd@NHNN&U8]fWPZdW:C[LH
>(LIUF2+)F?=?OA6b213HW[aQNM9+?8Z\(g+5P98#?XOCB(fa::JFe6c4FJ?_>=X
Q70g#YEL1O#b^?7?>fa+#-MLPD2SgS?b+>EZ:3=B831A,5ISEEGGLB@,Z[=:O@SQ
2EP&#F=UV7S>D=S9Bdd:?UX=W8[+3R=DbQ9ZgCPYSC1C&#,gU]<FVG8bZC9Ua:MZ
&<6]B:KF8I.6E/FODJKa4#SIR?7)E>\;SBf]?.N8<^@A>X;L@g4da2cA79#QWSAA
YdUVTL[g?HCUX3/-94U7bcPGQR0WP=L-X7.TH8(S(4_gKJ1ZF,^[LC0?\CCJ-WaJ
)20[1)&VJ8d=69Hd^b7^=fWc:RPAIU1M,V)9+2bDVV#^;;R<;a0f9A)^FG10##GB
d<XC0JV1XJICbdY>cI;VI?N.Z9W2LG&c9c0B[USTf^\?JB27X34]HHb,D0]11Y@b
ES6614[L7?U@;eN)Q\8DcG87,N(P;IE.6J_8c[Y]CZ^f<Lgb(6F0&N:]?9XLXZ1&
PH;AHS_gEL^M0[V?P4/,,/9C+ZgBXLCO_WI6LRSd5E&^ZWaX2ROJB8L[e&E@.F@&
F.]/cb#.5@?^UVY51KTJT1J2a3@Z7G_^E3CCARcD(KP:7(Qb\=](7)TL&7ET;JVe
^-6HWXP:HD?\GVH\+DW);2+&HQK76E5H-YWZDL5K;D/0=7G9D((4D;A<:f0W6@#Z
G^;?93g?@YKJA@2/FGdI]Gb07f&E\IeGD]Td;3NAV>Q>9Z5b@GYg@=K3>;(c&[BR
X#_QTe[0,D3(N_@d-ABD:UOgeQAgY]=Y.OUZ@UC/TC_Yf5O<F=FG8@bdS7B5_.(H
>SDc<OMGA[&Mg<^#EaXU0^+?,0S-^(W??8QHDcRd(19D_/]^3>Xa.:/>Q<OC)RTM
YJTEDcHT]/I:_3HS(_?UOe7;VQZW/>?;3c9;gOIEC)F]Td;06(ED;a5U@Y]Y#?Q+
.K_R=M?CZ:+;&7CIX-#d?QDaCe?O(KZDW-J9e9eS3B+LF>6f5O]W8Z1NOJ?T+HVS
?e1(3SV^O[8T7a#UE7GW/7^GL4)f3GF)e97WIb.O,V(O&RR/V?312^7(1<@cW<b3
6()TLWYXZX=I](d2ZB=>c=9Yd:gXA:bYe70D7<5H[gUV^fL?I]5/[KHAg1:Y<(?F
a3F-](\3Sc:/7HaHZ@-D#]PRQ#;?c=9a+0.N5aNcU>N-+T&fU;_>:3GbIAE5#76\
S:f8Q8G7PSA79Q81IBSKGYYC:5\BRa;N<aU9V0+A&06Ze,;>Ccf4JDU>WA&(Ge<E
YH=S,W#-[P<eR4.EE)6##0)BcL]g+N]eK[d6_L6OT4aQ)9IWb:D2>.U)AQL6)7R&
e5>Y+cLK/](>3O]BLDHZfV0/FF=UL(9GfOb_MC]EC59M0?H)XdF0R&X+#a9?_=OJ
TaO;&4f&E-)]:^EVL.C7]^7XR:QO2&V/G.LXS;Z]bd;]Dc\Te6BSb:DfJBZ-Q39S
DMWcb?2d:XScCeKF2Vd.eG#/9&<Y/<(AbMW>R\0(3=&Mf\[WA5=D6P#X9T?2R+?)
S9OYQ0A)P&KbX?8#9TMcADLJ1LH7NM09K5A#DSg:AJ5/BF:1B5SGD5O/]3.C7+@?
#f_<&@9>fIKO:RC./C#+6I.<M>V8)TZ,K0X3]B<.;YC<LeB=ZKWRV0,_2HDS-PW-
:XZ:UF#FAE@^\<<3;7>QX5?.M[NMT7^R2O_FXV-_09&,EKM9_>g2>(V/H<IC)3Ad
C?-65,0dIK@9&4?U:5DRQD:XD,UD,1QA>>CX+WQ^H8f^+C]Z#MQ=d52VU;TVX<DX
e[=LA(+HZ1Xgg/X,U7bD5a0e2_H(.C139>YNV4F,R2V&T&EKYLb)a<YA>c_6?D0P
4LJXV(LE\L_EG&aS>9:)3+E0DO87cg[B#UUP<]VJB5f6],ZO]:[XMDJ++,CVP=D+
NHGJT>2c:3Q10ZF??VH\A508-K,4]Zgab-#R]b_/;+LJGRM_bTWV(^fQE^SY1efR
6E1+VLIL/1T2&HTM10VFT9XTVgZJMSW(^S6MO5+R(G8fW.,]@PPe,F+Yf:A?K0TG
P-<63+\#+\W\5#K8#Q3F#+b+(6TRSc_/H)R0af5bgJ9)Jc+e6<,ASO,)/4Dag3_0
&g0+c6T4dG<BTaN@PS_OMZbZa:1&+dN-V(Y3K01K<TP2#d79L>?FXI3ef](P])0G
M5G5)..Q9-QQVZD&b7dFd3O^5J_cb.^X0eEH0&R,3LaO(CL1f)#9]bEA\(N7)6?Y
/AaFG],&PNZ]J(:IV)(GFg]UG1PVT5(R;$
`endprotected


